magic
tech gf180mcuD
magscale 1 5
timestamp 1702578009
<< obsm1 >>
rect 672 1538 9376 8262
<< metal2 >>
rect 2464 9600 2520 10000
rect 7392 9600 7448 10000
<< obsm2 >>
rect 854 9570 2434 9600
rect 2550 9570 7362 9600
rect 7478 9570 9362 9600
rect 854 625 9362 9570
<< metal3 >>
rect 0 9184 400 9240
rect 9600 8624 10000 8680
rect 0 7952 400 8008
rect 0 6720 400 6776
rect 9600 6160 10000 6216
rect 0 5488 400 5544
rect 0 4256 400 4312
rect 9600 3696 10000 3752
rect 0 3024 400 3080
rect 0 1792 400 1848
rect 9600 1232 10000 1288
rect 0 560 400 616
<< obsm3 >>
rect 430 9154 9600 9226
rect 400 8710 9600 9154
rect 400 8594 9570 8710
rect 400 8038 9600 8594
rect 430 7922 9600 8038
rect 400 6806 9600 7922
rect 430 6690 9600 6806
rect 400 6246 9600 6690
rect 400 6130 9570 6246
rect 400 5574 9600 6130
rect 430 5458 9600 5574
rect 400 4342 9600 5458
rect 430 4226 9600 4342
rect 400 3782 9600 4226
rect 400 3666 9570 3782
rect 400 3110 9600 3666
rect 430 2994 9600 3110
rect 400 1878 9600 2994
rect 430 1762 9600 1878
rect 400 1318 9600 1762
rect 400 1202 9570 1318
rect 400 646 9600 1202
rect 430 574 9600 646
<< metal4 >>
rect 1670 1538 1830 8262
rect 2748 1538 2908 8262
rect 3826 1538 3986 8262
rect 4904 1538 5064 8262
rect 5982 1538 6142 8262
rect 7060 1538 7220 8262
rect 8138 1538 8298 8262
rect 9216 1538 9376 8262
<< labels >>
rlabel metal2 s 2464 9600 2520 10000 6 clk
port 1 nsew signal input
rlabel metal2 s 7392 9600 7448 10000 6 reset
port 2 nsew signal input
rlabel metal3 s 0 3024 400 3080 6 rle1__input_r[0]
port 3 nsew signal input
rlabel metal3 s 0 4256 400 4312 6 rle1__input_r[1]
port 4 nsew signal input
rlabel metal3 s 0 5488 400 5544 6 rle1__input_r[2]
port 5 nsew signal input
rlabel metal3 s 0 6720 400 6776 6 rle1__input_r[3]
port 6 nsew signal input
rlabel metal3 s 0 7952 400 8008 6 rle1__input_r[4]
port 7 nsew signal input
rlabel metal3 s 0 9184 400 9240 6 rle1__input_r[5]
port 8 nsew signal input
rlabel metal3 s 0 560 400 616 6 rle1__input_r_rdy
port 9 nsew signal output
rlabel metal3 s 0 1792 400 1848 6 rle1__input_r_vld
port 10 nsew signal input
rlabel metal3 s 9600 6160 10000 6216 6 rle1__output_s[0]
port 11 nsew signal output
rlabel metal3 s 9600 8624 10000 8680 6 rle1__output_s[1]
port 12 nsew signal output
rlabel metal3 s 9600 1232 10000 1288 6 rle1__output_s_rdy
port 13 nsew signal input
rlabel metal3 s 9600 3696 10000 3752 6 rle1__output_s_vld
port 14 nsew signal output
rlabel metal4 s 1670 1538 1830 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 8262 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 8262 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 8262 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 8262 6 vss
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 368174
string GDS_FILE /home/proppy/src/github.com/proppy/xls-tapeouts/openlane/rle1_dec/runs/23_12_15_03_19/results/signoff/rle1_dec_wrap.magic.gds
string GDS_START 154096
<< end >>

