module __fmac__fmac_0_next(
  input wire clk,
  input wire reset,
  input wire [15:0] fmac__input_a,
  input wire fmac__input_a_vld,
  input wire [15:0] fmac__input_b,
  input wire fmac__input_b_vld,
  input wire fmac__reset,
  input wire fmac__reset_vld,
  input wire fmac__output_rdy,
  output wire [15:0] fmac__output,
  output wire fmac__output_vld,
  output wire fmac__input_a_rdy,
  output wire fmac__input_b_rdy,
  output wire fmac__reset_rdy
);
  // lint_off MULTIPLY
  function automatic [15:0] umul16b_8b_x_8b (input reg [7:0] lhs, input reg [7:0] rhs);
    begin
      umul16b_8b_x_8b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [15:0] __fmac__input_a_reg_init;
  assign __fmac__input_a_reg_init = {1'h0, 8'h00, 7'h00};
  wire [15:0] __fmac__input_b_reg_init;
  assign __fmac__input_b_reg_init = {1'h0, 8'h00, 7'h00};
  wire [15:0] __fmac__output_reg_init;
  assign __fmac__output_reg_init = {1'h0, 8'h00, 7'h00};
  reg [8:0] p0_result_exp__4;
  reg [15:0] p0_result_fraction__7;
  reg p0_result_sign__4;
  reg p0_literal_1952;
  reg p0_literal_1956;
  reg [7:0] p0_literal_1953;
  reg [6:0] ____state_2;
  reg [7:0] ____state_1;
  reg ____state_0;
  reg p0_valid;
  reg [15:0] __fmac__input_a_reg;
  reg __fmac__input_a_valid_reg;
  reg [15:0] __fmac__input_b_reg;
  reg __fmac__input_b_valid_reg;
  reg __fmac__reset_reg;
  reg __fmac__reset_valid_reg;
  reg [15:0] __fmac__output_reg;
  reg __fmac__output_valid_reg;
  wire [8:0] concat_2001;
  wire [7:0] wide_c__4;
  wire ugt_2005;
  wire [7:0] wide_c__3;
  wire [8:0] add_2009;
  wire [8:0] greater_exp;
  wire [8:0] add_2012;
  wire [24:0] wide_c__2;
  wire [8:0] sub_2014;
  wire [24:0] wide_ab;
  wire [8:0] sub_2016;
  wire [8:0] rshift_c;
  wire [24:0] dropped_c;
  wire [24:0] dropped_ab;
  wire [7:0] dropped_c__2;
  wire [8:0] rshift_ab;
  wire [24:0] shifted_ab;
  wire [24:0] sticky_ab;
  wire [24:0] shifted_c;
  wire [24:0] sticky_c;
  wire [24:0] or_2037;
  wire [24:0] or_2039;
  wire greater_sign;
  wire [25:0] neg_2045;
  wire [25:0] neg_2047;
  wire [26:0] shifted_ab__1;
  wire [26:0] shifted_c__1;
  wire [26:0] shifted_ab__2;
  wire [26:0] shifted_c__2;
  wire [26:0] sum_fraction;
  wire [25:0] abs_fraction__1;
  wire [25:0] reverse_2061;
  wire [26:0] one_hot_2062;
  wire [4:0] encode_2063;
  wire __stateancel__2;
  wire __statearry_bit;
  wire [25:0] leading_zeroes;
  wire [24:0] __statearry_fraction__2;
  wire [25:0] add_2080;
  wire [2:0] concat_2081;
  wire [24:0] __statearry_fraction__1;
  wire [24:0] __stateancel_fraction;
  wire [24:0] shifted_fraction;
  wire [16:0] normal_chunk;
  wire [16:0] half_of_extra;
  wire [1:0] half_way_chunk;
  wire [8:0] concat_2093;
  wire do_round_up;
  wire [8:0] add_2096;
  wire [8:0] rounded_fraction__1;
  wire [6:0] a_fraction__3;
  wire [7:0] a_bexp__4;
  wire [6:0] b_fraction__3;
  wire [7:0] b_bexp__4;
  wire rounding_carry;
  wire [7:0] a_fraction__4;
  wire [7:0] b_fraction__4;
  wire [9:0] add_2103;
  wire [7:0] a_fraction__5;
  wire [7:0] b_fraction__5;
  wire [9:0] add_2107;
  wire [15:0] fraction;
  wire [9:0] bexp__4;
  wire [9:0] bexp__5;
  wire [8:0] add_1907;
  wire eq_1910;
  wire eq_1911;
  wire [8:0] high_exp__2;
  wire [9:0] bexp__11;
  wire [9:0] bexp__12;
  wire eq_2116;
  wire eq_2117;
  wire [7:0] max_exp__8;
  wire [7:0] max_exp__6;
  wire [9:0] bexp__13;
  wire ne_2125;
  wire and_2126;
  wire eq_2127;
  wire eq_2128;
  wire [9:0] bexp__14;
  wire p1_all_active_states_valid;
  wire [8:0] bexp__6;
  wire [7:0] max_exp;
  wire [7:0] max_exp__5;
  wire p1_stage_valid;
  wire fmac__output_valid_inv;
  wire has_pos_inf;
  wire has_neg_inf;
  wire fraction_is_zero;
  wire eq_1921;
  wire eq_1923;
  wire __fmac__output_vld_buf;
  wire fmac__output_valid_load_en;
  wire and_2148;
  wire and_reduce_2153;
  wire and_1929;
  wire and_1930;
  wire [8:0] result_exp__3;
  wire fmac__output_load_en;
  wire p1_all_active_states_ready;
  wire is_result_nan__2;
  wire is_operand_inf;
  wire result_sign__1;
  wire has_0_arg;
  wire has_inf_arg;
  wire [15:0] fraction__1;
  wire [8:0] sub_exp;
  wire p1_stage_done;
  wire p1_not_valid;
  wire p0_all_active_states_valid;
  wire p0_all_active_inputs_valid;
  wire p0_all_active_outputs_ready;
  wire p0_all_active_states_ready;
  wire result_sign__2;
  wire [6:0] result_fraction__1;
  wire is_subnormal;
  wire p0_enable;
  wire p0_stage_done;
  wire result_sign__5;
  wire [7:0] max_exp__7;
  wire [6:0] result_fraction__3;
  wire is_result_nan__1;
  wire [15:0] result_fraction__5;
  wire a_sign__2;
  wire b_sign__2;
  wire p0_data_enable;
  wire fmac__input_a_valid_inv;
  wire fmac__input_b_valid_inv;
  wire fmac__reset_valid_inv;
  wire [7:0] result_exp__2;
  wire [6:0] result_fraction__4;
  wire [8:0] high_exp;
  wire [15:0] result_fraction__6;
  wire [15:0] nan_fraction;
  wire result_sign__3;
  wire fmac__input_a_valid_load_en;
  wire fmac__input_b_valid_load_en;
  wire fmac__reset_valid_load_en;
  wire nor_2184;
  wire [7:0] and_2186;
  wire [6:0] and_2188;
  wire [8:0] result_exp__4;
  wire [15:0] result_fraction__7;
  wire result_sign__4;
  wire literal_1952;
  wire literal_1956;
  wire [7:0] literal_1953;
  wire fmac__input_a_load_en;
  wire fmac__input_b_load_en;
  wire fmac__reset_load_en;
  wire [15:0] acc__1;
  assign concat_2001 = {p0_literal_1956, ____state_1};
  assign wide_c__4 = {p0_literal_1952, ____state_2} | 8'h80;
  assign ugt_2005 = p0_result_exp__4 > concat_2001;
  assign wide_c__3 = wide_c__4 & {8{____state_1 != p0_literal_1953}};
  assign add_2009 = concat_2001 + 9'h019;
  assign greater_exp = ugt_2005 ? p0_result_exp__4 : concat_2001;
  assign add_2012 = p0_result_exp__4 + 9'h019;
  assign wide_c__2 = {wide_c__3, 17'h0_0000};
  assign sub_2014 = add_2009 - greater_exp;
  assign wide_ab = {p0_result_fraction__7, 9'h000};
  assign sub_2016 = add_2012 - greater_exp;
  assign rshift_c = greater_exp - concat_2001;
  assign dropped_c = sub_2014 >= 9'h019 ? 25'h000_0000 : wide_c__2 << sub_2014;
  assign dropped_ab = sub_2016 >= 9'h019 ? 25'h000_0000 : wide_ab << sub_2016;
  assign dropped_c__2 = rshift_c > 9'h018 ? wide_c__3 : dropped_c[24:17];
  assign rshift_ab = greater_exp - p0_result_exp__4;
  assign shifted_ab = rshift_ab >= 9'h019 ? 25'h000_0000 : wide_ab >> rshift_ab;
  assign sticky_ab = {24'h00_0000, dropped_ab[24:9] != 16'h0000};
  assign shifted_c = rshift_c >= 9'h019 ? 25'h000_0000 : wide_c__2 >> rshift_c;
  assign sticky_c = {24'h00_0000, dropped_c__2 != 8'h00};
  assign or_2037 = shifted_ab | sticky_ab;
  assign or_2039 = shifted_c | sticky_c;
  assign greater_sign = ugt_2005 ? p0_result_sign__4 : ____state_0;
  assign neg_2045 = -{1'h0, or_2037};
  assign neg_2047 = -{1'h0, or_2039};
  assign shifted_ab__1 = {2'h0, or_2037};
  assign shifted_c__1 = {2'h0, or_2039};
  assign shifted_ab__2 = p0_result_sign__4 ^ greater_sign ? {{1{neg_2045[25]}}, neg_2045} : shifted_ab__1;
  assign shifted_c__2 = ____state_0 ^ greater_sign ? {{1{neg_2047[25]}}, neg_2047} : shifted_c__1;
  assign sum_fraction = shifted_ab__2 + shifted_c__2;
  assign abs_fraction__1 = sum_fraction[26] ? -sum_fraction[25:0] : sum_fraction[25:0];
  assign reverse_2061 = {abs_fraction__1[0], abs_fraction__1[1], abs_fraction__1[2], abs_fraction__1[3], abs_fraction__1[4], abs_fraction__1[5], abs_fraction__1[6], abs_fraction__1[7], abs_fraction__1[8], abs_fraction__1[9], abs_fraction__1[10], abs_fraction__1[11], abs_fraction__1[12], abs_fraction__1[13], abs_fraction__1[14], abs_fraction__1[15], abs_fraction__1[16], abs_fraction__1[17], abs_fraction__1[18], abs_fraction__1[19], abs_fraction__1[20], abs_fraction__1[21], abs_fraction__1[22], abs_fraction__1[23], abs_fraction__1[24], abs_fraction__1[25]};
  assign one_hot_2062 = {reverse_2061[25:0] == 26'h000_0000, reverse_2061[25] && reverse_2061[24:0] == 25'h000_0000, reverse_2061[24] && reverse_2061[23:0] == 24'h00_0000, reverse_2061[23] && reverse_2061[22:0] == 23'h00_0000, reverse_2061[22] && reverse_2061[21:0] == 22'h00_0000, reverse_2061[21] && reverse_2061[20:0] == 21'h00_0000, reverse_2061[20] && reverse_2061[19:0] == 20'h0_0000, reverse_2061[19] && reverse_2061[18:0] == 19'h0_0000, reverse_2061[18] && reverse_2061[17:0] == 18'h0_0000, reverse_2061[17] && reverse_2061[16:0] == 17'h0_0000, reverse_2061[16] && reverse_2061[15:0] == 16'h0000, reverse_2061[15] && reverse_2061[14:0] == 15'h0000, reverse_2061[14] && reverse_2061[13:0] == 14'h0000, reverse_2061[13] && reverse_2061[12:0] == 13'h0000, reverse_2061[12] && reverse_2061[11:0] == 12'h000, reverse_2061[11] && reverse_2061[10:0] == 11'h000, reverse_2061[10] && reverse_2061[9:0] == 10'h000, reverse_2061[9] && reverse_2061[8:0] == 9'h000, reverse_2061[8] && reverse_2061[7:0] == 8'h00, reverse_2061[7] && reverse_2061[6:0] == 7'h00, reverse_2061[6] && reverse_2061[5:0] == 6'h00, reverse_2061[5] && reverse_2061[4:0] == 5'h00, reverse_2061[4] && reverse_2061[3:0] == 4'h0, reverse_2061[3] && reverse_2061[2:0] == 3'h0, reverse_2061[2] && reverse_2061[1:0] == 2'h0, reverse_2061[1] && !reverse_2061[0], reverse_2061[0]};
  assign encode_2063 = {one_hot_2062[16] | one_hot_2062[17] | one_hot_2062[18] | one_hot_2062[19] | one_hot_2062[20] | one_hot_2062[21] | one_hot_2062[22] | one_hot_2062[23] | one_hot_2062[24] | one_hot_2062[25] | one_hot_2062[26], one_hot_2062[8] | one_hot_2062[9] | one_hot_2062[10] | one_hot_2062[11] | one_hot_2062[12] | one_hot_2062[13] | one_hot_2062[14] | one_hot_2062[15] | one_hot_2062[24] | one_hot_2062[25] | one_hot_2062[26], one_hot_2062[4] | one_hot_2062[5] | one_hot_2062[6] | one_hot_2062[7] | one_hot_2062[12] | one_hot_2062[13] | one_hot_2062[14] | one_hot_2062[15] | one_hot_2062[20] | one_hot_2062[21] | one_hot_2062[22] | one_hot_2062[23], one_hot_2062[2] | one_hot_2062[3] | one_hot_2062[6] | one_hot_2062[7] | one_hot_2062[10] | one_hot_2062[11] | one_hot_2062[14] | one_hot_2062[15] | one_hot_2062[18] | one_hot_2062[19] | one_hot_2062[22] | one_hot_2062[23] | one_hot_2062[26], one_hot_2062[1] | one_hot_2062[3] | one_hot_2062[5] | one_hot_2062[7] | one_hot_2062[9] | one_hot_2062[11] | one_hot_2062[13] | one_hot_2062[15] | one_hot_2062[17] | one_hot_2062[19] | one_hot_2062[21] | one_hot_2062[23] | one_hot_2062[25]};
  assign __stateancel__2 = |encode_2063[4:1];
  assign __statearry_bit = abs_fraction__1[25];
  assign leading_zeroes = {21'h00_0000, encode_2063};
  assign __statearry_fraction__2 = abs_fraction__1[25:1];
  assign add_2080 = leading_zeroes + 26'h3ff_ffff;
  assign concat_2081 = {~(__statearry_bit | __stateancel__2), ~(__statearry_bit | ~__stateancel__2), ~(~__statearry_bit | __stateancel__2)};
  assign __statearry_fraction__1 = __statearry_fraction__2 | {24'h00_0000, abs_fraction__1[0]};
  assign __stateancel_fraction = add_2080 >= 26'h000_0019 ? 25'h000_0000 : abs_fraction__1[24:0] << add_2080;
  assign shifted_fraction = __statearry_fraction__1 & {25{concat_2081[0]}} | __stateancel_fraction & {25{concat_2081[1]}} | abs_fraction__1[24:0] & {25{concat_2081[2]}};
  assign normal_chunk = shifted_fraction[16:0];
  assign half_of_extra = 17'h1_0000;
  assign half_way_chunk = shifted_fraction[17:16];
  assign concat_2093 = {1'h0, shifted_fraction[24:17]};
  assign do_round_up = normal_chunk > half_of_extra | half_way_chunk == 2'h3;
  assign add_2096 = concat_2093 + 9'h001;
  assign rounded_fraction__1 = do_round_up ? add_2096 : concat_2093;
  assign a_fraction__3 = __fmac__input_a_reg[6:0];
  assign a_bexp__4 = __fmac__input_a_reg[14:7];
  assign b_fraction__3 = __fmac__input_b_reg[6:0];
  assign b_bexp__4 = __fmac__input_b_reg[14:7];
  assign rounding_carry = rounded_fraction__1[8];
  assign a_fraction__4 = {1'h0, a_fraction__3} | 8'h80;
  assign b_fraction__4 = {1'h0, b_fraction__3} | 8'h80;
  assign add_2103 = {1'h0, greater_exp} + {9'h000, rounding_carry};
  assign a_fraction__5 = a_fraction__4 & {8{a_bexp__4 != 8'h00}};
  assign b_fraction__5 = b_fraction__4 & {8{b_bexp__4 != 8'h00}};
  assign add_2107 = add_2103 + 10'h001;
  assign fraction = umul16b_8b_x_8b(a_fraction__5, b_fraction__5);
  assign bexp__4 = add_2107 - {5'h00, encode_2063};
  assign bexp__5 = bexp__4 & {10{sum_fraction != 27'h000_0000}};
  assign add_1907 = {1'h0, a_bexp__4} + {1'h0, b_bexp__4};
  assign eq_1910 = a_bexp__4 == 8'h00;
  assign eq_1911 = b_bexp__4 == 8'h00;
  assign high_exp__2 = 9'h1ff;
  assign bexp__11 = {1'h0, add_1907};
  assign bexp__12 = {9'h000, fraction[15]} + 10'h381;
  assign eq_2116 = p0_result_exp__4 == high_exp__2;
  assign eq_2117 = p0_result_fraction__7 == 16'h0000;
  assign max_exp__8 = 8'hff;
  assign max_exp__6 = 8'hff;
  assign bexp__13 = bexp__11 + bexp__12;
  assign ne_2125 = ____state_2 != 7'h00;
  assign and_2126 = eq_2116 & eq_2117;
  assign eq_2127 = ____state_1 == max_exp__6;
  assign eq_2128 = ____state_2 == 7'h00;
  assign bexp__14 = bexp__13 & {10{~(eq_1910 | eq_1911)}};
  assign p1_all_active_states_valid = 1'h1;
  assign bexp__6 = bexp__5[8:0] & {9{~bexp__5[9]}};
  assign max_exp = 8'hff;
  assign max_exp__5 = 8'hff;
  assign p1_stage_valid = p1_all_active_states_valid & p0_valid;
  assign fmac__output_valid_inv = ~__fmac__output_valid_reg;
  assign has_pos_inf = ~(~(eq_2116 & eq_2117) | p0_result_sign__4) | ~(____state_1 != max_exp__8 | ne_2125 | ____state_0);
  assign has_neg_inf = and_2126 & p0_result_sign__4 | eq_2127 & eq_2128 & ____state_0;
  assign fraction_is_zero = sum_fraction == 27'h000_0000;
  assign eq_1921 = a_bexp__4 == max_exp;
  assign eq_1923 = b_bexp__4 == max_exp__5;
  assign __fmac__output_vld_buf = __fmac__reset_valid_reg & p1_stage_valid & 1'h1;
  assign fmac__output_valid_load_en = fmac__output_rdy | fmac__output_valid_inv;
  assign and_2148 = eq_2127 & eq_2128;
  assign and_reduce_2153 = &bexp__6[7:0];
  assign and_1929 = eq_1921 & a_fraction__3 == 7'h00;
  assign and_1930 = eq_1923 & b_fraction__3 == 7'h00;
  assign result_exp__3 = bexp__14[8:0] & {9{$signed(bexp__14) > $signed(10'h000)}};
  assign fmac__output_load_en = __fmac__output_vld_buf & fmac__output_valid_load_en;
  assign p1_all_active_states_ready = 1'h1;
  assign is_result_nan__2 = eq_2116 & p0_result_fraction__7 != 16'h0000 | eq_2127 & ne_2125 | has_pos_inf & has_neg_inf;
  assign is_operand_inf = and_2126 | and_2148;
  assign result_sign__1 = ~(~sum_fraction[26] | greater_sign) | ~(sum_fraction[26] | fraction_is_zero | ~greater_sign);
  assign has_0_arg = eq_1910 | eq_1911;
  assign has_inf_arg = and_1929 | and_1930;
  assign fraction__1 = fraction[15] ? fraction : {fraction[14:0], 1'h0};
  assign sub_exp = bexp__14[9] ? -bexp__14[8:0] : bexp__14[8:0];
  assign p1_stage_done = p1_stage_valid & __fmac__reset_valid_reg & fmac__output_load_en & p1_all_active_states_ready;
  assign p1_not_valid = ~p0_valid;
  assign p0_all_active_states_valid = 1'h1;
  assign p0_all_active_inputs_valid = __fmac__input_a_valid_reg & __fmac__input_b_valid_reg;
  assign p0_all_active_outputs_ready = 1'h1;
  assign p0_all_active_states_ready = 1'h1;
  assign result_sign__2 = is_operand_inf ? ~has_pos_inf : result_sign__1;
  assign result_fraction__1 = rounded_fraction__1[6:0];
  assign is_subnormal = $signed(bexp__14) <= $signed(10'h000);
  assign p0_enable = p1_stage_done | p1_not_valid;
  assign p0_stage_done = p0_all_active_states_valid & p0_all_active_inputs_valid & p0_all_active_outputs_ready & p0_all_active_states_ready;
  assign result_sign__5 = ~is_result_nan__2 & result_sign__2;
  assign max_exp__7 = 8'hff;
  assign result_fraction__3 = result_fraction__1 & {7{bexp__6 != 9'h000}} & {7{~(bexp__6[8] | and_reduce_2153)}} & {7{~(and_2126 | and_2148)}};
  assign is_result_nan__1 = eq_1921 & a_fraction__3 != 7'h00 | eq_1923 & b_fraction__3 != 7'h00 | has_0_arg & has_inf_arg;
  assign result_fraction__5 = is_subnormal ? (sub_exp >= 9'h010 ? 16'h0000 : fraction__1 >> sub_exp) : fraction__1;
  assign a_sign__2 = __fmac__input_a_reg[15:15];
  assign b_sign__2 = __fmac__input_b_reg[15:15];
  assign p0_data_enable = p0_enable & p0_stage_done;
  assign fmac__input_a_valid_inv = ~__fmac__input_a_valid_reg;
  assign fmac__input_b_valid_inv = ~__fmac__input_b_valid_reg;
  assign fmac__reset_valid_inv = ~__fmac__reset_valid_reg;
  assign result_exp__2 = is_result_nan__2 | is_operand_inf | bexp__6[8] | and_reduce_2153 ? max_exp__7 : bexp__6[7:0];
  assign result_fraction__4 = is_result_nan__2 ? 7'h08 : result_fraction__3;
  assign high_exp = 9'h1ff;
  assign result_fraction__6 = result_fraction__5 & {16{~(&result_exp__3)}} & {16{~(and_1929 | and_1930)}};
  assign nan_fraction = 16'h0001;
  assign result_sign__3 = a_sign__2 ^ b_sign__2;
  assign fmac__input_a_valid_load_en = p0_data_enable | fmac__input_a_valid_inv;
  assign fmac__input_b_valid_load_en = p0_data_enable | fmac__input_b_valid_inv;
  assign fmac__reset_valid_load_en = p1_stage_done | fmac__reset_valid_inv;
  assign nor_2184 = ~(__fmac__reset_reg | ~result_sign__5);
  assign and_2186 = result_exp__2 & {8{~__fmac__reset_reg}};
  assign and_2188 = result_fraction__4 & {7{~__fmac__reset_reg}};
  assign result_exp__4 = is_result_nan__1 | has_inf_arg ? high_exp : result_exp__3;
  assign result_fraction__7 = is_result_nan__1 ? nan_fraction : result_fraction__6;
  assign result_sign__4 = ~is_result_nan__1 & result_sign__3;
  assign literal_1952 = 1'h0;
  assign literal_1956 = 1'h0;
  assign literal_1953 = 8'h00;
  assign fmac__input_a_load_en = fmac__input_a_vld & fmac__input_a_valid_load_en;
  assign fmac__input_b_load_en = fmac__input_b_vld & fmac__input_b_valid_load_en;
  assign fmac__reset_load_en = fmac__reset_vld & fmac__reset_valid_load_en;
  assign acc__1 = {nor_2184, and_2186, and_2188};
  always_ff @ (posedge clk) begin
    if (reset) begin
      p0_result_exp__4 <= 9'h000;
      p0_result_fraction__7 <= 16'h0000;
      p0_result_sign__4 <= 1'h0;
      p0_literal_1952 <= 1'h0;
      p0_literal_1956 <= 1'h0;
      p0_literal_1953 <= 8'h00;
      ____state_2 <= 7'h00;
      ____state_1 <= 8'h00;
      ____state_0 <= 1'h0;
      p0_valid <= 1'h0;
      __fmac__input_a_reg <= __fmac__input_a_reg_init;
      __fmac__input_a_valid_reg <= 1'h0;
      __fmac__input_b_reg <= __fmac__input_b_reg_init;
      __fmac__input_b_valid_reg <= 1'h0;
      __fmac__reset_reg <= 1'h0;
      __fmac__reset_valid_reg <= 1'h0;
      __fmac__output_reg <= __fmac__output_reg_init;
      __fmac__output_valid_reg <= 1'h0;
    end else begin
      p0_result_exp__4 <= p0_data_enable ? result_exp__4 : p0_result_exp__4;
      p0_result_fraction__7 <= p0_data_enable ? result_fraction__7 : p0_result_fraction__7;
      p0_result_sign__4 <= p0_data_enable ? result_sign__4 : p0_result_sign__4;
      p0_literal_1952 <= p0_data_enable ? literal_1952 : p0_literal_1952;
      p0_literal_1956 <= p0_data_enable ? literal_1956 : p0_literal_1956;
      p0_literal_1953 <= p0_data_enable ? literal_1953 : p0_literal_1953;
      ____state_2 <= p1_stage_done ? and_2188 : ____state_2;
      ____state_1 <= p1_stage_done ? and_2186 : ____state_1;
      ____state_0 <= p1_stage_done ? nor_2184 : ____state_0;
      p0_valid <= p0_enable ? p0_stage_done : p0_valid;
      __fmac__input_a_reg <= fmac__input_a_load_en ? fmac__input_a : __fmac__input_a_reg;
      __fmac__input_a_valid_reg <= fmac__input_a_valid_load_en ? fmac__input_a_vld : __fmac__input_a_valid_reg;
      __fmac__input_b_reg <= fmac__input_b_load_en ? fmac__input_b : __fmac__input_b_reg;
      __fmac__input_b_valid_reg <= fmac__input_b_valid_load_en ? fmac__input_b_vld : __fmac__input_b_valid_reg;
      __fmac__reset_reg <= fmac__reset_load_en ? fmac__reset : __fmac__reset_reg;
      __fmac__reset_valid_reg <= fmac__reset_valid_load_en ? fmac__reset_vld : __fmac__reset_valid_reg;
      __fmac__output_reg <= fmac__output_load_en ? acc__1 : __fmac__output_reg;
      __fmac__output_valid_reg <= fmac__output_valid_load_en ? __fmac__output_vld_buf : __fmac__output_valid_reg;
    end
  end
  carry_and_cancel: assert property (@(posedge clk) disable iff (reset) ~p1_stage_done | ~(__statearry_bit & __stateancel__2)) else $fatal(0, "Assertion failure via fail! @ /home/proppy/xls-env/share/xls/xls/dslx/ir_convert/ir_converter_main.runfiles/com_google_xls/xls/dslx/stdlib/apfloat.x:2152:15-2152:56");
  assign fmac__output = __fmac__output_reg;
  assign fmac__output_vld = __fmac__output_valid_reg;
  assign fmac__input_a_rdy = fmac__input_a_load_en;
  assign fmac__input_b_rdy = fmac__input_b_load_en;
  assign fmac__reset_rdy = fmac__reset_load_en;
endmodule
