magic
tech gf180mcuD
magscale 1 10
timestamp 1702516874
<< obsm1 >>
rect 1344 3076 58731 26850
<< metal2 >>
rect 9856 29200 9968 30000
rect 29792 29200 29904 30000
rect 49728 29200 49840 30000
<< obsm2 >>
rect 1260 29140 9796 29200
rect 10028 29140 29732 29200
rect 29964 29140 49668 29200
rect 49900 29140 58703 29200
rect 1260 1362 58703 29140
<< metal3 >>
rect 0 28224 800 28336
rect 59200 27328 60000 27440
rect 0 26432 800 26544
rect 0 24640 800 24752
rect 59200 23744 60000 23856
rect 0 22848 800 22960
rect 0 21056 800 21168
rect 59200 20160 60000 20272
rect 0 19264 800 19376
rect 0 17472 800 17584
rect 59200 16576 60000 16688
rect 0 15680 800 15792
rect 0 13888 800 14000
rect 59200 12992 60000 13104
rect 0 12096 800 12208
rect 0 10304 800 10416
rect 59200 9408 60000 9520
rect 0 8512 800 8624
rect 0 6720 800 6832
rect 59200 5824 60000 5936
rect 0 4928 800 5040
rect 0 3136 800 3248
rect 59200 2240 60000 2352
rect 0 1344 800 1456
<< obsm3 >>
rect 860 28164 59332 28308
rect 800 27500 59332 28164
rect 800 27268 59140 27500
rect 800 26604 59332 27268
rect 860 26372 59332 26604
rect 800 24812 59332 26372
rect 860 24580 59332 24812
rect 800 23916 59332 24580
rect 800 23684 59140 23916
rect 800 23020 59332 23684
rect 860 22788 59332 23020
rect 800 21228 59332 22788
rect 860 20996 59332 21228
rect 800 20332 59332 20996
rect 800 20100 59140 20332
rect 800 19436 59332 20100
rect 860 19204 59332 19436
rect 800 17644 59332 19204
rect 860 17412 59332 17644
rect 800 16748 59332 17412
rect 800 16516 59140 16748
rect 800 15852 59332 16516
rect 860 15620 59332 15852
rect 800 14060 59332 15620
rect 860 13828 59332 14060
rect 800 13164 59332 13828
rect 800 12932 59140 13164
rect 800 12268 59332 12932
rect 860 12036 59332 12268
rect 800 10476 59332 12036
rect 860 10244 59332 10476
rect 800 9580 59332 10244
rect 800 9348 59140 9580
rect 800 8684 59332 9348
rect 860 8452 59332 8684
rect 800 6892 59332 8452
rect 860 6660 59332 6892
rect 800 5996 59332 6660
rect 800 5764 59140 5996
rect 800 5100 59332 5764
rect 860 4868 59332 5100
rect 800 3308 59332 4868
rect 860 3076 59332 3308
rect 800 2412 59332 3076
rect 800 2180 59140 2412
rect 800 1516 59332 2180
rect 860 1372 59332 1516
<< metal4 >>
rect 8337 3076 8657 26716
rect 15490 3076 15810 26716
rect 22644 3076 22964 26716
rect 29797 3076 30117 26716
rect 36951 3076 37271 26716
rect 44104 3076 44424 26716
rect 51258 3076 51578 26716
rect 58411 3076 58731 26716
<< obsm4 >>
rect 1820 5394 8277 26302
rect 8717 5394 15430 26302
rect 15870 5394 22584 26302
rect 23024 5394 29737 26302
rect 30177 5394 36891 26302
rect 37331 5394 44044 26302
rect 44484 5394 51198 26302
rect 51638 5394 55972 26302
<< labels >>
rlabel metal3 s 0 1344 800 1456 6 a[0]
port 1 nsew signal input
rlabel metal3 s 0 3136 800 3248 6 a[1]
port 2 nsew signal input
rlabel metal3 s 0 4928 800 5040 6 a[2]
port 3 nsew signal input
rlabel metal3 s 0 6720 800 6832 6 a[3]
port 4 nsew signal input
rlabel metal3 s 0 8512 800 8624 6 a[4]
port 5 nsew signal input
rlabel metal3 s 0 10304 800 10416 6 a[5]
port 6 nsew signal input
rlabel metal3 s 0 12096 800 12208 6 a[6]
port 7 nsew signal input
rlabel metal3 s 0 13888 800 14000 6 a[7]
port 8 nsew signal input
rlabel metal3 s 0 15680 800 15792 6 b[0]
port 9 nsew signal input
rlabel metal3 s 0 17472 800 17584 6 b[1]
port 10 nsew signal input
rlabel metal3 s 0 19264 800 19376 6 b[2]
port 11 nsew signal input
rlabel metal3 s 0 21056 800 21168 6 b[3]
port 12 nsew signal input
rlabel metal3 s 0 22848 800 22960 6 b[4]
port 13 nsew signal input
rlabel metal3 s 0 24640 800 24752 6 b[5]
port 14 nsew signal input
rlabel metal3 s 0 26432 800 26544 6 b[6]
port 15 nsew signal input
rlabel metal3 s 0 28224 800 28336 6 b[7]
port 16 nsew signal input
rlabel metal2 s 9856 29200 9968 30000 6 op[0]
port 17 nsew signal input
rlabel metal2 s 29792 29200 29904 30000 6 op[1]
port 18 nsew signal input
rlabel metal2 s 49728 29200 49840 30000 6 op[2]
port 19 nsew signal input
rlabel metal3 s 59200 2240 60000 2352 6 out[0]
port 20 nsew signal output
rlabel metal3 s 59200 5824 60000 5936 6 out[1]
port 21 nsew signal output
rlabel metal3 s 59200 9408 60000 9520 6 out[2]
port 22 nsew signal output
rlabel metal3 s 59200 12992 60000 13104 6 out[3]
port 23 nsew signal output
rlabel metal3 s 59200 16576 60000 16688 6 out[4]
port 24 nsew signal output
rlabel metal3 s 59200 20160 60000 20272 6 out[5]
port 25 nsew signal output
rlabel metal3 s 59200 23744 60000 23856 6 out[6]
port 26 nsew signal output
rlabel metal3 s 59200 27328 60000 27440 6 out[7]
port 27 nsew signal output
rlabel metal4 s 8337 3076 8657 26716 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 22644 3076 22964 26716 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 36951 3076 37271 26716 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 51258 3076 51578 26716 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 15490 3076 15810 26716 6 vss
port 29 nsew ground bidirectional
rlabel metal4 s 29797 3076 30117 26716 6 vss
port 29 nsew ground bidirectional
rlabel metal4 s 44104 3076 44424 26716 6 vss
port 29 nsew ground bidirectional
rlabel metal4 s 58411 3076 58731 26716 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1769250
string GDS_FILE /home/proppy/src/github.com/proppy/xls-tapeouts/openlane/fpu8/runs/23_12_14_10_19/results/signoff/fpu8_wrap.magic.gds
string GDS_START 451064
<< end >>

