magic
tech gf180mcuD
magscale 1 5
timestamp 1702516938
<< obsm1 >>
rect 672 1538 9376 8262
<< metal2 >>
rect 2464 9600 2520 10000
rect 7392 9600 7448 10000
<< obsm2 >>
rect 854 9570 2434 9600
rect 2550 9570 7362 9600
rect 7478 9570 9362 9600
rect 854 569 9362 9570
<< metal3 >>
rect 9600 9184 10000 9240
rect 0 8624 400 8680
rect 9600 7952 10000 8008
rect 9600 6720 10000 6776
rect 0 6160 400 6216
rect 9600 5488 10000 5544
rect 9600 4256 10000 4312
rect 0 3696 400 3752
rect 9600 3024 10000 3080
rect 9600 1792 10000 1848
rect 0 1232 400 1288
rect 9600 560 10000 616
<< obsm3 >>
rect 400 9154 9570 9226
rect 400 8710 9600 9154
rect 430 8594 9600 8710
rect 400 8038 9600 8594
rect 400 7922 9570 8038
rect 400 6806 9600 7922
rect 400 6690 9570 6806
rect 400 6246 9600 6690
rect 430 6130 9600 6246
rect 400 5574 9600 6130
rect 400 5458 9570 5574
rect 400 4342 9600 5458
rect 400 4226 9570 4342
rect 400 3782 9600 4226
rect 430 3666 9600 3782
rect 400 3110 9600 3666
rect 400 2994 9570 3110
rect 400 1878 9600 2994
rect 400 1762 9570 1878
rect 400 1318 9600 1762
rect 430 1202 9600 1318
rect 400 646 9600 1202
rect 400 574 9570 646
<< metal4 >>
rect 1670 1538 1830 8262
rect 2748 1538 2908 8262
rect 3826 1538 3986 8262
rect 4904 1538 5064 8262
rect 5982 1538 6142 8262
rect 7060 1538 7220 8262
rect 8138 1538 8298 8262
rect 9216 1538 9376 8262
<< obsm4 >>
rect 2982 2529 3796 7047
rect 4016 2529 4874 7047
rect 5094 2529 5922 7047
<< labels >>
rlabel metal2 s 2464 9600 2520 10000 6 clk
port 1 nsew signal input
rlabel metal2 s 7392 9600 7448 10000 6 reset
port 2 nsew signal input
rlabel metal3 s 0 6160 400 6216 6 rle1__input_r[0]
port 3 nsew signal input
rlabel metal3 s 0 8624 400 8680 6 rle1__input_r[1]
port 4 nsew signal input
rlabel metal3 s 0 1232 400 1288 6 rle1__input_r_rdy
port 5 nsew signal output
rlabel metal3 s 0 3696 400 3752 6 rle1__input_r_vld
port 6 nsew signal input
rlabel metal3 s 9600 3024 10000 3080 6 rle1__output_s[0]
port 7 nsew signal output
rlabel metal3 s 9600 4256 10000 4312 6 rle1__output_s[1]
port 8 nsew signal output
rlabel metal3 s 9600 5488 10000 5544 6 rle1__output_s[2]
port 9 nsew signal output
rlabel metal3 s 9600 6720 10000 6776 6 rle1__output_s[3]
port 10 nsew signal output
rlabel metal3 s 9600 7952 10000 8008 6 rle1__output_s[4]
port 11 nsew signal output
rlabel metal3 s 9600 9184 10000 9240 6 rle1__output_s[5]
port 12 nsew signal output
rlabel metal3 s 9600 560 10000 616 6 rle1__output_s_rdy
port 13 nsew signal input
rlabel metal3 s 9600 1792 10000 1848 6 rle1__output_s_vld
port 14 nsew signal output
rlabel metal4 s 1670 1538 1830 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 8262 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 8262 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 8262 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 8262 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 8262 6 vss
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 411060
string GDS_FILE /home/proppy/src/github.com/proppy/xls-tapeouts/openlane/rle1_enc/runs/23_12_14_10_21/results/signoff/rle1_enc_wrap.magic.gds
string GDS_START 174002
<< end >>

