magic
tech gf180mcuD
magscale 1 5
timestamp 1702578008
<< metal1 >>
rect 672 8245 9296 8262
rect 672 8219 1685 8245
rect 1711 8219 1737 8245
rect 1763 8219 1789 8245
rect 1815 8219 3841 8245
rect 3867 8219 3893 8245
rect 3919 8219 3945 8245
rect 3971 8219 5997 8245
rect 6023 8219 6049 8245
rect 6075 8219 6101 8245
rect 6127 8219 8153 8245
rect 8179 8219 8205 8245
rect 8231 8219 8257 8245
rect 8283 8219 9296 8245
rect 672 8202 9296 8219
rect 7457 8135 7463 8161
rect 7489 8135 7495 8161
rect 1191 8049 1217 8055
rect 8073 8023 8079 8049
rect 8105 8023 8111 8049
rect 8577 8023 8583 8049
rect 8609 8023 8615 8049
rect 1191 8017 1217 8023
rect 855 7993 881 7999
rect 855 7961 881 7967
rect 1583 7993 1609 7999
rect 1583 7961 1609 7967
rect 1023 7937 1049 7943
rect 1023 7905 1049 7911
rect 1359 7937 1385 7943
rect 1359 7905 1385 7911
rect 8471 7937 8497 7943
rect 8471 7905 8497 7911
rect 672 7853 9376 7870
rect 672 7827 2763 7853
rect 2789 7827 2815 7853
rect 2841 7827 2867 7853
rect 2893 7827 4919 7853
rect 4945 7827 4971 7853
rect 4997 7827 5023 7853
rect 5049 7827 7075 7853
rect 7101 7827 7127 7853
rect 7153 7827 7179 7853
rect 7205 7827 9231 7853
rect 9257 7827 9283 7853
rect 9309 7827 9335 7853
rect 9361 7827 9376 7853
rect 672 7810 9376 7827
rect 1079 7769 1105 7775
rect 1079 7737 1105 7743
rect 8359 7769 8385 7775
rect 8359 7737 8385 7743
rect 1415 7713 1441 7719
rect 1415 7681 1441 7687
rect 1471 7657 1497 7663
rect 2865 7631 2871 7657
rect 2897 7631 2903 7657
rect 6393 7631 6399 7657
rect 6425 7631 6431 7657
rect 6617 7631 6623 7657
rect 6649 7631 6655 7657
rect 1471 7625 1497 7631
rect 3201 7575 3207 7601
rect 3233 7575 3239 7601
rect 4265 7575 4271 7601
rect 4297 7575 4303 7601
rect 4937 7575 4943 7601
rect 4969 7575 4975 7601
rect 6001 7575 6007 7601
rect 6033 7575 6039 7601
rect 7009 7575 7015 7601
rect 7041 7575 7047 7601
rect 8073 7575 8079 7601
rect 8105 7575 8111 7601
rect 672 7461 9296 7478
rect 672 7435 1685 7461
rect 1711 7435 1737 7461
rect 1763 7435 1789 7461
rect 1815 7435 3841 7461
rect 3867 7435 3893 7461
rect 3919 7435 3945 7461
rect 3971 7435 5997 7461
rect 6023 7435 6049 7461
rect 6075 7435 6101 7461
rect 6127 7435 8153 7461
rect 8179 7435 8205 7461
rect 8231 7435 8257 7461
rect 8283 7435 9296 7461
rect 672 7418 9296 7435
rect 1415 7321 1441 7327
rect 1415 7289 1441 7295
rect 3599 7321 3625 7327
rect 7295 7321 7321 7327
rect 5553 7295 5559 7321
rect 5585 7295 5591 7321
rect 3599 7289 3625 7295
rect 7295 7289 7321 7295
rect 3263 7265 3289 7271
rect 3655 7265 3681 7271
rect 6063 7265 6089 7271
rect 3145 7239 3151 7265
rect 3177 7239 3183 7265
rect 3425 7239 3431 7265
rect 3457 7239 3463 7265
rect 3761 7239 3767 7265
rect 3793 7239 3799 7265
rect 4097 7239 4103 7265
rect 4129 7239 4135 7265
rect 3263 7233 3289 7239
rect 3655 7233 3681 7239
rect 6063 7233 6089 7239
rect 6959 7265 6985 7271
rect 6959 7233 6985 7239
rect 7071 7265 7097 7271
rect 7071 7233 7097 7239
rect 7239 7265 7265 7271
rect 7239 7233 7265 7239
rect 3039 7209 3065 7215
rect 5727 7209 5753 7215
rect 4489 7183 4495 7209
rect 4521 7183 4527 7209
rect 3039 7177 3065 7183
rect 5727 7177 5753 7183
rect 5839 7209 5865 7215
rect 5839 7177 5865 7183
rect 7351 7209 7377 7215
rect 7351 7177 7377 7183
rect 7463 7209 7489 7215
rect 7463 7177 7489 7183
rect 7575 7209 7601 7215
rect 7575 7177 7601 7183
rect 7631 7209 7657 7215
rect 7631 7177 7657 7183
rect 1471 7153 1497 7159
rect 5895 7153 5921 7159
rect 3201 7127 3207 7153
rect 3233 7127 3239 7153
rect 1471 7121 1497 7127
rect 5895 7121 5921 7127
rect 672 7069 9376 7086
rect 672 7043 2763 7069
rect 2789 7043 2815 7069
rect 2841 7043 2867 7069
rect 2893 7043 4919 7069
rect 4945 7043 4971 7069
rect 4997 7043 5023 7069
rect 5049 7043 7075 7069
rect 7101 7043 7127 7069
rect 7153 7043 7179 7069
rect 7205 7043 9231 7069
rect 9257 7043 9283 7069
rect 9309 7043 9335 7069
rect 9361 7043 9376 7069
rect 672 7026 9376 7043
rect 5111 6985 5137 6991
rect 3313 6959 3319 6985
rect 3345 6959 3351 6985
rect 5111 6953 5137 6959
rect 5447 6985 5473 6991
rect 5447 6953 5473 6959
rect 5727 6985 5753 6991
rect 5727 6953 5753 6959
rect 5839 6985 5865 6991
rect 5839 6953 5865 6959
rect 7071 6985 7097 6991
rect 7071 6953 7097 6959
rect 1023 6929 1049 6935
rect 1023 6897 1049 6903
rect 1471 6929 1497 6935
rect 1471 6897 1497 6903
rect 2479 6929 2505 6935
rect 2479 6897 2505 6903
rect 2647 6929 2673 6935
rect 2647 6897 2673 6903
rect 2983 6929 3009 6935
rect 5223 6929 5249 6935
rect 3649 6903 3655 6929
rect 3681 6903 3687 6929
rect 3985 6903 3991 6929
rect 4017 6903 4023 6929
rect 2983 6897 3009 6903
rect 5223 6897 5249 6903
rect 5559 6929 5585 6935
rect 5559 6897 5585 6903
rect 5615 6929 5641 6935
rect 6959 6929 6985 6935
rect 6169 6903 6175 6929
rect 6201 6903 6207 6929
rect 5615 6897 5641 6903
rect 6959 6897 6985 6903
rect 855 6873 881 6879
rect 4999 6873 5025 6879
rect 2865 6847 2871 6873
rect 2897 6847 2903 6873
rect 3201 6847 3207 6873
rect 3233 6847 3239 6873
rect 3537 6847 3543 6873
rect 3569 6847 3575 6873
rect 3873 6847 3879 6873
rect 3905 6847 3911 6873
rect 855 6841 881 6847
rect 4999 6841 5025 6847
rect 5335 6873 5361 6879
rect 5335 6841 5361 6847
rect 5895 6873 5921 6879
rect 6511 6873 6537 6879
rect 6113 6847 6119 6873
rect 6145 6847 6151 6873
rect 5895 6841 5921 6847
rect 6511 6841 6537 6847
rect 6679 6873 6705 6879
rect 6679 6841 6705 6847
rect 6903 6873 6929 6879
rect 6903 6841 6929 6847
rect 1247 6817 1273 6823
rect 1247 6785 1273 6791
rect 1415 6761 1441 6767
rect 1415 6729 1441 6735
rect 672 6677 9296 6694
rect 672 6651 1685 6677
rect 1711 6651 1737 6677
rect 1763 6651 1789 6677
rect 1815 6651 3841 6677
rect 3867 6651 3893 6677
rect 3919 6651 3945 6677
rect 3971 6651 5997 6677
rect 6023 6651 6049 6677
rect 6075 6651 6101 6677
rect 6127 6651 8153 6677
rect 8179 6651 8205 6677
rect 8231 6651 8257 6677
rect 8283 6651 9296 6677
rect 672 6634 9296 6651
rect 5447 6593 5473 6599
rect 5447 6561 5473 6567
rect 6791 6593 6817 6599
rect 6791 6561 6817 6567
rect 8975 6537 9001 6543
rect 2529 6511 2535 6537
rect 2561 6511 2567 6537
rect 8975 6505 9001 6511
rect 7463 6481 7489 6487
rect 1129 6455 1135 6481
rect 1161 6455 1167 6481
rect 4545 6455 4551 6481
rect 4577 6455 4583 6481
rect 5161 6455 5167 6481
rect 5193 6455 5199 6481
rect 6729 6455 6735 6481
rect 6761 6455 6767 6481
rect 7569 6455 7575 6481
rect 7601 6455 7607 6481
rect 8017 6455 8023 6481
rect 8049 6455 8055 6481
rect 7463 6449 7489 6455
rect 5615 6425 5641 6431
rect 1465 6399 1471 6425
rect 1497 6399 1503 6425
rect 5049 6399 5055 6425
rect 5081 6399 5087 6425
rect 5615 6393 5641 6399
rect 5839 6425 5865 6431
rect 5839 6393 5865 6399
rect 7239 6425 7265 6431
rect 7345 6399 7351 6425
rect 7377 6399 7383 6425
rect 7239 6393 7265 6399
rect 6007 6369 6033 6375
rect 4657 6343 4663 6369
rect 4689 6343 4695 6369
rect 6007 6337 6033 6343
rect 6847 6369 6873 6375
rect 6847 6337 6873 6343
rect 6959 6369 6985 6375
rect 7457 6343 7463 6369
rect 7489 6343 7495 6369
rect 6959 6337 6985 6343
rect 672 6285 9376 6302
rect 672 6259 2763 6285
rect 2789 6259 2815 6285
rect 2841 6259 2867 6285
rect 2893 6259 4919 6285
rect 4945 6259 4971 6285
rect 4997 6259 5023 6285
rect 5049 6259 7075 6285
rect 7101 6259 7127 6285
rect 7153 6259 7179 6285
rect 7205 6259 9231 6285
rect 9257 6259 9283 6285
rect 9309 6259 9335 6285
rect 9361 6259 9376 6285
rect 672 6242 9376 6259
rect 1639 6201 1665 6207
rect 1639 6169 1665 6175
rect 4495 6201 4521 6207
rect 4495 6169 4521 6175
rect 4775 6201 4801 6207
rect 4775 6169 4801 6175
rect 4831 6201 4857 6207
rect 4831 6169 4857 6175
rect 6623 6201 6649 6207
rect 6623 6169 6649 6175
rect 6903 6201 6929 6207
rect 7687 6201 7713 6207
rect 7233 6175 7239 6201
rect 7265 6175 7271 6201
rect 6903 6169 6929 6175
rect 7687 6169 7713 6175
rect 7967 6201 7993 6207
rect 7967 6169 7993 6175
rect 6007 6145 6033 6151
rect 1297 6119 1303 6145
rect 1329 6119 1335 6145
rect 1689 6119 1695 6145
rect 1721 6119 1727 6145
rect 5217 6119 5223 6145
rect 5249 6119 5255 6145
rect 6007 6113 6033 6119
rect 6119 6145 6145 6151
rect 6119 6113 6145 6119
rect 6343 6145 6369 6151
rect 6343 6113 6369 6119
rect 8023 6145 8049 6151
rect 8023 6113 8049 6119
rect 1415 6089 1441 6095
rect 1073 6063 1079 6089
rect 1105 6063 1111 6089
rect 1415 6057 1441 6063
rect 1583 6089 1609 6095
rect 2255 6089 2281 6095
rect 3319 6089 3345 6095
rect 5111 6089 5137 6095
rect 6063 6089 6089 6095
rect 6847 6089 6873 6095
rect 1969 6063 1975 6089
rect 2001 6063 2007 6089
rect 2361 6063 2367 6089
rect 2393 6063 2399 6089
rect 3481 6063 3487 6089
rect 3513 6063 3519 6089
rect 4265 6063 4271 6089
rect 4297 6063 4303 6089
rect 4377 6063 4383 6089
rect 4409 6063 4415 6089
rect 4937 6063 4943 6089
rect 4969 6063 4975 6089
rect 5329 6063 5335 6089
rect 5361 6063 5367 6089
rect 5609 6063 5615 6089
rect 5641 6063 5647 6089
rect 5833 6063 5839 6089
rect 5865 6063 5871 6089
rect 6225 6063 6231 6089
rect 6257 6063 6263 6089
rect 1583 6057 1609 6063
rect 2255 6057 2281 6063
rect 3319 6057 3345 6063
rect 5111 6057 5137 6063
rect 6063 6057 6089 6063
rect 6847 6057 6873 6063
rect 7407 6089 7433 6095
rect 7407 6057 7433 6063
rect 1359 6033 1385 6039
rect 1359 6001 1385 6007
rect 3375 6033 3401 6039
rect 3375 6001 3401 6007
rect 1191 5977 1217 5983
rect 2199 5977 2225 5983
rect 1857 5951 1863 5977
rect 1889 5951 1895 5977
rect 1191 5945 1217 5951
rect 2199 5945 2225 5951
rect 4551 5977 4577 5983
rect 4551 5945 4577 5951
rect 6511 5977 6537 5983
rect 6511 5945 6537 5951
rect 6679 5977 6705 5983
rect 6679 5945 6705 5951
rect 6903 5977 6929 5983
rect 6903 5945 6929 5951
rect 7575 5977 7601 5983
rect 7575 5945 7601 5951
rect 7743 5977 7769 5983
rect 7743 5945 7769 5951
rect 7911 5977 7937 5983
rect 7911 5945 7937 5951
rect 672 5893 9296 5910
rect 672 5867 1685 5893
rect 1711 5867 1737 5893
rect 1763 5867 1789 5893
rect 1815 5867 3841 5893
rect 3867 5867 3893 5893
rect 3919 5867 3945 5893
rect 3971 5867 5997 5893
rect 6023 5867 6049 5893
rect 6075 5867 6101 5893
rect 6127 5867 8153 5893
rect 8179 5867 8205 5893
rect 8231 5867 8257 5893
rect 8283 5867 9296 5893
rect 672 5850 9296 5867
rect 6175 5753 6201 5759
rect 1465 5727 1471 5753
rect 1497 5727 1503 5753
rect 2529 5727 2535 5753
rect 2561 5727 2567 5753
rect 4097 5727 4103 5753
rect 4129 5727 4135 5753
rect 9081 5727 9087 5753
rect 9113 5727 9119 5753
rect 6175 5721 6201 5727
rect 6287 5697 6313 5703
rect 1129 5671 1135 5697
rect 1161 5671 1167 5697
rect 5833 5671 5839 5697
rect 5865 5671 5871 5697
rect 6841 5671 6847 5697
rect 6873 5671 6879 5697
rect 7625 5671 7631 5697
rect 7657 5671 7663 5697
rect 6287 5665 6313 5671
rect 6735 5641 6761 5647
rect 6735 5609 6761 5615
rect 6959 5641 6985 5647
rect 6959 5609 6985 5615
rect 7127 5641 7153 5647
rect 8017 5615 8023 5641
rect 8049 5615 8055 5641
rect 7127 5609 7153 5615
rect 7015 5585 7041 5591
rect 6449 5559 6455 5585
rect 6481 5559 6487 5585
rect 7015 5553 7041 5559
rect 7183 5585 7209 5591
rect 7183 5553 7209 5559
rect 7239 5585 7265 5591
rect 7239 5553 7265 5559
rect 672 5501 9376 5518
rect 672 5475 2763 5501
rect 2789 5475 2815 5501
rect 2841 5475 2867 5501
rect 2893 5475 4919 5501
rect 4945 5475 4971 5501
rect 4997 5475 5023 5501
rect 5049 5475 7075 5501
rect 7101 5475 7127 5501
rect 7153 5475 7179 5501
rect 7205 5475 9231 5501
rect 9257 5475 9283 5501
rect 9309 5475 9335 5501
rect 9361 5475 9376 5501
rect 672 5458 9376 5475
rect 1247 5417 1273 5423
rect 1247 5385 1273 5391
rect 4495 5417 4521 5423
rect 4495 5385 4521 5391
rect 4887 5417 4913 5423
rect 8129 5391 8135 5417
rect 8161 5391 8167 5417
rect 4887 5385 4913 5391
rect 855 5361 881 5367
rect 855 5329 881 5335
rect 1023 5361 1049 5367
rect 1023 5329 1049 5335
rect 2199 5361 2225 5367
rect 2199 5329 2225 5335
rect 2311 5361 2337 5367
rect 2311 5329 2337 5335
rect 2647 5361 2673 5367
rect 2647 5329 2673 5335
rect 4999 5361 5025 5367
rect 6169 5335 6175 5361
rect 6201 5335 6207 5361
rect 4999 5329 5025 5335
rect 4719 5305 4745 5311
rect 7911 5305 7937 5311
rect 8415 5305 8441 5311
rect 2473 5279 2479 5305
rect 2505 5279 2511 5305
rect 2809 5279 2815 5305
rect 2841 5279 2847 5305
rect 5161 5279 5167 5305
rect 5193 5279 5199 5305
rect 8073 5279 8079 5305
rect 8105 5279 8111 5305
rect 4719 5273 4745 5279
rect 7911 5273 7937 5279
rect 8415 5273 8441 5279
rect 8695 5305 8721 5311
rect 8695 5273 8721 5279
rect 1415 5249 1441 5255
rect 4831 5249 4857 5255
rect 2137 5223 2143 5249
rect 2169 5223 2175 5249
rect 3201 5223 3207 5249
rect 3233 5223 3239 5249
rect 4265 5223 4271 5249
rect 4297 5223 4303 5249
rect 1415 5217 1441 5223
rect 4831 5217 4857 5223
rect 8303 5249 8329 5255
rect 8303 5217 8329 5223
rect 8751 5249 8777 5255
rect 8751 5217 8777 5223
rect 8975 5249 9001 5255
rect 8975 5217 9001 5223
rect 1471 5193 1497 5199
rect 1471 5161 1497 5167
rect 2479 5193 2505 5199
rect 2479 5161 2505 5167
rect 8191 5193 8217 5199
rect 8191 5161 8217 5167
rect 8919 5193 8945 5199
rect 8919 5161 8945 5167
rect 672 5109 9296 5126
rect 672 5083 1685 5109
rect 1711 5083 1737 5109
rect 1763 5083 1789 5109
rect 1815 5083 3841 5109
rect 3867 5083 3893 5109
rect 3919 5083 3945 5109
rect 3971 5083 5997 5109
rect 6023 5083 6049 5109
rect 6075 5083 6101 5109
rect 6127 5083 8153 5109
rect 8179 5083 8205 5109
rect 8231 5083 8257 5109
rect 8283 5083 9296 5109
rect 672 5066 9296 5083
rect 7127 5025 7153 5031
rect 3201 4999 3207 5025
rect 3233 4999 3239 5025
rect 7127 4993 7153 4999
rect 3543 4969 3569 4975
rect 6399 4969 6425 4975
rect 2529 4943 2535 4969
rect 2561 4943 2567 4969
rect 4881 4943 4887 4969
rect 4913 4943 4919 4969
rect 5609 4943 5615 4969
rect 5641 4943 5647 4969
rect 3543 4937 3569 4943
rect 6399 4937 6425 4943
rect 7239 4969 7265 4975
rect 7905 4943 7911 4969
rect 7937 4943 7943 4969
rect 9025 4943 9031 4969
rect 9057 4943 9063 4969
rect 7239 4937 7265 4943
rect 6287 4913 6313 4919
rect 1129 4887 1135 4913
rect 1161 4887 1167 4913
rect 3257 4887 3263 4913
rect 3289 4887 3295 4913
rect 4433 4887 4439 4913
rect 4465 4887 4471 4913
rect 4825 4887 4831 4913
rect 4857 4887 4863 4913
rect 5273 4887 5279 4913
rect 5305 4887 5311 4913
rect 5441 4887 5447 4913
rect 5473 4887 5479 4913
rect 6001 4887 6007 4913
rect 6033 4887 6039 4913
rect 6287 4881 6313 4887
rect 6511 4913 6537 4919
rect 7351 4913 7377 4919
rect 6897 4887 6903 4913
rect 6929 4887 6935 4913
rect 7009 4887 7015 4913
rect 7041 4887 7047 4913
rect 7569 4887 7575 4913
rect 7601 4887 7607 4913
rect 6511 4881 6537 4887
rect 7351 4881 7377 4887
rect 2927 4857 2953 4863
rect 6175 4857 6201 4863
rect 1465 4831 1471 4857
rect 1497 4831 1503 4857
rect 3033 4831 3039 4857
rect 3065 4831 3071 4857
rect 4209 4831 4215 4857
rect 4241 4831 4247 4857
rect 4769 4831 4775 4857
rect 4801 4831 4807 4857
rect 5497 4831 5503 4857
rect 5529 4831 5535 4857
rect 2927 4825 2953 4831
rect 6175 4825 6201 4831
rect 4047 4801 4073 4807
rect 7407 4801 7433 4807
rect 3089 4775 3095 4801
rect 3121 4775 3127 4801
rect 4545 4775 4551 4801
rect 4577 4775 4583 4801
rect 4047 4769 4073 4775
rect 7407 4769 7433 4775
rect 672 4717 9376 4734
rect 672 4691 2763 4717
rect 2789 4691 2815 4717
rect 2841 4691 2867 4717
rect 2893 4691 4919 4717
rect 4945 4691 4971 4717
rect 4997 4691 5023 4717
rect 5049 4691 7075 4717
rect 7101 4691 7127 4717
rect 7153 4691 7179 4717
rect 7205 4691 9231 4717
rect 9257 4691 9283 4717
rect 9309 4691 9335 4717
rect 9361 4691 9376 4717
rect 672 4674 9376 4691
rect 1471 4633 1497 4639
rect 1471 4601 1497 4607
rect 4383 4633 4409 4639
rect 4383 4601 4409 4607
rect 4887 4633 4913 4639
rect 4887 4601 4913 4607
rect 1023 4577 1049 4583
rect 1023 4545 1049 4551
rect 1863 4577 1889 4583
rect 1863 4545 1889 4551
rect 2031 4577 2057 4583
rect 2031 4545 2057 4551
rect 2815 4577 2841 4583
rect 2815 4545 2841 4551
rect 2983 4577 3009 4583
rect 2983 4545 3009 4551
rect 3151 4577 3177 4583
rect 3151 4545 3177 4551
rect 4495 4577 4521 4583
rect 4495 4545 4521 4551
rect 5559 4577 5585 4583
rect 8751 4577 8777 4583
rect 7569 4551 7575 4577
rect 7601 4551 7607 4577
rect 5559 4545 5585 4551
rect 8751 4545 8777 4551
rect 855 4521 881 4527
rect 1695 4521 1721 4527
rect 4271 4521 4297 4527
rect 1465 4495 1471 4521
rect 1497 4495 1503 4521
rect 2137 4495 2143 4521
rect 2169 4495 2175 4521
rect 2361 4495 2367 4521
rect 2393 4495 2399 4521
rect 3313 4495 3319 4521
rect 3345 4495 3351 4521
rect 855 4489 881 4495
rect 1695 4489 1721 4495
rect 4271 4489 4297 4495
rect 4327 4521 4353 4527
rect 4327 4489 4353 4495
rect 4831 4521 4857 4527
rect 4831 4489 4857 4495
rect 4943 4521 4969 4527
rect 4943 4489 4969 4495
rect 5111 4521 5137 4527
rect 5111 4489 5137 4495
rect 5223 4521 5249 4527
rect 5223 4489 5249 4495
rect 5447 4521 5473 4527
rect 8695 4521 8721 4527
rect 6225 4495 6231 4521
rect 6257 4495 6263 4521
rect 5447 4489 5473 4495
rect 8695 4489 8721 4495
rect 8863 4521 8889 4527
rect 8863 4489 8889 4495
rect 1247 4465 1273 4471
rect 1247 4433 1273 4439
rect 2087 4465 2113 4471
rect 2087 4433 2113 4439
rect 3207 4465 3233 4471
rect 3207 4433 3233 4439
rect 5335 4465 5361 4471
rect 5335 4433 5361 4439
rect 1639 4409 1665 4415
rect 2305 4383 2311 4409
rect 2337 4383 2343 4409
rect 1639 4377 1665 4383
rect 672 4325 9296 4342
rect 672 4299 1685 4325
rect 1711 4299 1737 4325
rect 1763 4299 1789 4325
rect 1815 4299 3841 4325
rect 3867 4299 3893 4325
rect 3919 4299 3945 4325
rect 3971 4299 5997 4325
rect 6023 4299 6049 4325
rect 6075 4299 6101 4325
rect 6127 4299 8153 4325
rect 8179 4299 8205 4325
rect 8231 4299 8257 4325
rect 8283 4299 9296 4325
rect 672 4282 9296 4299
rect 5447 4241 5473 4247
rect 5447 4209 5473 4215
rect 6903 4241 6929 4247
rect 6903 4209 6929 4215
rect 1465 4159 1471 4185
rect 1497 4159 1503 4185
rect 2529 4159 2535 4185
rect 2561 4159 2567 4185
rect 3817 4159 3823 4185
rect 3849 4159 3855 4185
rect 4881 4159 4887 4185
rect 4913 4159 4919 4185
rect 5049 4159 5055 4185
rect 5081 4159 5087 4185
rect 6785 4159 6791 4185
rect 6817 4159 6823 4185
rect 7849 4159 7855 4185
rect 7881 4159 7887 4185
rect 8913 4159 8919 4185
rect 8945 4159 8951 4185
rect 5335 4129 5361 4135
rect 1129 4103 1135 4129
rect 1161 4103 1167 4129
rect 3425 4103 3431 4129
rect 3457 4103 3463 4129
rect 5335 4097 5361 4103
rect 5559 4129 5585 4135
rect 5559 4097 5585 4103
rect 5783 4129 5809 4135
rect 5783 4097 5809 4103
rect 6231 4129 6257 4135
rect 6231 4097 6257 4103
rect 6343 4129 6369 4135
rect 6449 4103 6455 4129
rect 6481 4103 6487 4129
rect 7513 4103 7519 4129
rect 7545 4103 7551 4129
rect 6343 4097 6369 4103
rect 5671 4073 5697 4079
rect 5671 4041 5697 4047
rect 5895 4073 5921 4079
rect 5895 4041 5921 4047
rect 5951 4073 5977 4079
rect 7065 4047 7071 4073
rect 7097 4047 7103 4073
rect 5951 4041 5977 4047
rect 6175 4017 6201 4023
rect 6175 3985 6201 3991
rect 6287 4017 6313 4023
rect 6287 3985 6313 3991
rect 6791 4017 6817 4023
rect 6791 3985 6817 3991
rect 7239 4017 7265 4023
rect 7239 3985 7265 3991
rect 672 3933 9376 3950
rect 672 3907 2763 3933
rect 2789 3907 2815 3933
rect 2841 3907 2867 3933
rect 2893 3907 4919 3933
rect 4945 3907 4971 3933
rect 4997 3907 5023 3933
rect 5049 3907 7075 3933
rect 7101 3907 7127 3933
rect 7153 3907 7179 3933
rect 7205 3907 9231 3933
rect 9257 3907 9283 3933
rect 9309 3907 9335 3933
rect 9361 3907 9376 3933
rect 672 3890 9376 3907
rect 1471 3849 1497 3855
rect 1471 3817 1497 3823
rect 2703 3849 2729 3855
rect 4495 3849 4521 3855
rect 3369 3823 3375 3849
rect 3401 3823 3407 3849
rect 5105 3823 5111 3849
rect 5137 3823 5143 3849
rect 2703 3817 2729 3823
rect 4495 3817 4521 3823
rect 1415 3793 1441 3799
rect 4719 3793 4745 3799
rect 3761 3767 3767 3793
rect 3793 3767 3799 3793
rect 1415 3761 1441 3767
rect 4719 3761 4745 3767
rect 4831 3793 4857 3799
rect 4831 3761 4857 3767
rect 5335 3793 5361 3799
rect 5335 3761 5361 3767
rect 6623 3793 6649 3799
rect 6623 3761 6649 3767
rect 8863 3793 8889 3799
rect 8863 3761 8889 3767
rect 2927 3737 2953 3743
rect 2927 3705 2953 3711
rect 2983 3737 3009 3743
rect 2983 3705 3009 3711
rect 3207 3737 3233 3743
rect 4215 3737 4241 3743
rect 3313 3711 3319 3737
rect 3345 3711 3351 3737
rect 3873 3711 3879 3737
rect 3905 3711 3911 3737
rect 3207 3705 3233 3711
rect 4215 3705 4241 3711
rect 4887 3737 4913 3743
rect 8639 3737 8665 3743
rect 5049 3711 5055 3737
rect 5081 3711 5087 3737
rect 6953 3711 6959 3737
rect 6985 3711 6991 3737
rect 7345 3711 7351 3737
rect 7377 3711 7383 3737
rect 4887 3705 4913 3711
rect 8639 3705 8665 3711
rect 8975 3737 9001 3743
rect 8975 3705 9001 3711
rect 2423 3681 2449 3687
rect 2423 3649 2449 3655
rect 3095 3681 3121 3687
rect 3095 3649 3121 3655
rect 8303 3681 8329 3687
rect 8303 3649 8329 3655
rect 8751 3681 8777 3687
rect 8751 3649 8777 3655
rect 672 3541 9296 3558
rect 672 3515 1685 3541
rect 1711 3515 1737 3541
rect 1763 3515 1789 3541
rect 1815 3515 3841 3541
rect 3867 3515 3893 3541
rect 3919 3515 3945 3541
rect 3971 3515 5997 3541
rect 6023 3515 6049 3541
rect 6075 3515 6101 3541
rect 6127 3515 8153 3541
rect 8179 3515 8205 3541
rect 8231 3515 8257 3541
rect 8283 3515 9296 3541
rect 672 3498 9296 3515
rect 4937 3431 4943 3457
rect 4969 3431 4975 3457
rect 6225 3431 6231 3457
rect 6257 3431 6263 3457
rect 6791 3401 6817 3407
rect 3201 3375 3207 3401
rect 3233 3375 3239 3401
rect 4265 3375 4271 3401
rect 4297 3375 4303 3401
rect 5833 3375 5839 3401
rect 5865 3375 5871 3401
rect 6791 3369 6817 3375
rect 8975 3401 9001 3407
rect 8975 3369 9001 3375
rect 1415 3345 1441 3351
rect 1415 3313 1441 3319
rect 1471 3345 1497 3351
rect 6399 3345 6425 3351
rect 2865 3319 2871 3345
rect 2897 3319 2903 3345
rect 4545 3319 4551 3345
rect 4577 3319 4583 3345
rect 4993 3319 4999 3345
rect 5025 3319 5031 3345
rect 5217 3319 5223 3345
rect 5249 3319 5255 3345
rect 5777 3319 5783 3345
rect 5809 3319 5815 3345
rect 6169 3319 6175 3345
rect 6201 3319 6207 3345
rect 7177 3319 7183 3345
rect 7209 3319 7215 3345
rect 7513 3319 7519 3345
rect 7545 3319 7551 3345
rect 7905 3319 7911 3345
rect 7937 3319 7943 3345
rect 1471 3313 1497 3319
rect 6399 3313 6425 3319
rect 855 3289 881 3295
rect 855 3257 881 3263
rect 1023 3289 1049 3295
rect 1023 3257 1049 3263
rect 6735 3289 6761 3295
rect 6735 3257 6761 3263
rect 6847 3289 6873 3295
rect 7065 3263 7071 3289
rect 7097 3263 7103 3289
rect 6847 3257 6873 3263
rect 1247 3233 1273 3239
rect 1247 3201 1273 3207
rect 672 3149 9376 3166
rect 672 3123 2763 3149
rect 2789 3123 2815 3149
rect 2841 3123 2867 3149
rect 2893 3123 4919 3149
rect 4945 3123 4971 3149
rect 4997 3123 5023 3149
rect 5049 3123 7075 3149
rect 7101 3123 7127 3149
rect 7153 3123 7179 3149
rect 7205 3123 9231 3149
rect 9257 3123 9283 3149
rect 9309 3123 9335 3149
rect 9361 3123 9376 3149
rect 672 3106 9376 3123
rect 7183 3065 7209 3071
rect 7183 3033 7209 3039
rect 7463 3065 7489 3071
rect 8751 3065 8777 3071
rect 7737 3039 7743 3065
rect 7769 3039 7775 3065
rect 7463 3033 7489 3039
rect 8751 3033 8777 3039
rect 6505 2983 6511 3009
rect 6537 2983 6543 3009
rect 8129 2983 8135 3009
rect 8161 2983 8167 3009
rect 6897 2927 6903 2953
rect 6929 2927 6935 2953
rect 7737 2927 7743 2953
rect 7769 2927 7775 2953
rect 8185 2927 8191 2953
rect 8217 2927 8223 2953
rect 5447 2897 5473 2903
rect 5447 2865 5473 2871
rect 7071 2897 7097 2903
rect 7407 2897 7433 2903
rect 7177 2871 7183 2897
rect 7209 2871 7215 2897
rect 7071 2865 7097 2871
rect 7407 2865 7433 2871
rect 672 2757 9296 2774
rect 672 2731 1685 2757
rect 1711 2731 1737 2757
rect 1763 2731 1789 2757
rect 1815 2731 3841 2757
rect 3867 2731 3893 2757
rect 3919 2731 3945 2757
rect 3971 2731 5997 2757
rect 6023 2731 6049 2757
rect 6075 2731 6101 2757
rect 6127 2731 8153 2757
rect 8179 2731 8205 2757
rect 8231 2731 8257 2757
rect 8283 2731 9296 2757
rect 672 2714 9296 2731
rect 2983 2673 3009 2679
rect 2983 2641 3009 2647
rect 7295 2673 7321 2679
rect 7295 2641 7321 2647
rect 6847 2617 6873 2623
rect 6847 2585 6873 2591
rect 2927 2561 2953 2567
rect 2927 2529 2953 2535
rect 7351 2561 7377 2567
rect 7351 2529 7377 2535
rect 672 2365 9376 2382
rect 672 2339 2763 2365
rect 2789 2339 2815 2365
rect 2841 2339 2867 2365
rect 2893 2339 4919 2365
rect 4945 2339 4971 2365
rect 4997 2339 5023 2365
rect 5049 2339 7075 2365
rect 7101 2339 7127 2365
rect 7153 2339 7179 2365
rect 7205 2339 9231 2365
rect 9257 2339 9283 2365
rect 9309 2339 9335 2365
rect 9361 2339 9376 2365
rect 672 2322 9376 2339
rect 1023 2281 1049 2287
rect 1023 2249 1049 2255
rect 855 2169 881 2175
rect 855 2137 881 2143
rect 1247 2113 1273 2119
rect 1247 2081 1273 2087
rect 672 1973 9296 1990
rect 672 1947 1685 1973
rect 1711 1947 1737 1973
rect 1763 1947 1789 1973
rect 1815 1947 3841 1973
rect 3867 1947 3893 1973
rect 3919 1947 3945 1973
rect 3971 1947 5997 1973
rect 6023 1947 6049 1973
rect 6075 1947 6101 1973
rect 6127 1947 8153 1973
rect 8179 1947 8205 1973
rect 8231 1947 8257 1973
rect 8283 1947 9296 1973
rect 672 1930 9296 1947
rect 967 1833 993 1839
rect 967 1801 993 1807
rect 2137 1751 2143 1777
rect 2169 1751 2175 1777
rect 8807 1721 8833 1727
rect 9087 1721 9113 1727
rect 8913 1695 8919 1721
rect 8945 1695 8951 1721
rect 8807 1689 8833 1695
rect 9087 1689 9113 1695
rect 672 1581 9376 1598
rect 672 1555 2763 1581
rect 2789 1555 2815 1581
rect 2841 1555 2867 1581
rect 2893 1555 4919 1581
rect 4945 1555 4971 1581
rect 4997 1555 5023 1581
rect 5049 1555 7075 1581
rect 7101 1555 7127 1581
rect 7153 1555 7179 1581
rect 7205 1555 9231 1581
rect 9257 1555 9283 1581
rect 9309 1555 9335 1581
rect 9361 1555 9376 1581
rect 672 1538 9376 1555
<< via1 >>
rect 1685 8219 1711 8245
rect 1737 8219 1763 8245
rect 1789 8219 1815 8245
rect 3841 8219 3867 8245
rect 3893 8219 3919 8245
rect 3945 8219 3971 8245
rect 5997 8219 6023 8245
rect 6049 8219 6075 8245
rect 6101 8219 6127 8245
rect 8153 8219 8179 8245
rect 8205 8219 8231 8245
rect 8257 8219 8283 8245
rect 7463 8135 7489 8161
rect 1191 8023 1217 8049
rect 8079 8023 8105 8049
rect 8583 8023 8609 8049
rect 855 7967 881 7993
rect 1583 7967 1609 7993
rect 1023 7911 1049 7937
rect 1359 7911 1385 7937
rect 8471 7911 8497 7937
rect 2763 7827 2789 7853
rect 2815 7827 2841 7853
rect 2867 7827 2893 7853
rect 4919 7827 4945 7853
rect 4971 7827 4997 7853
rect 5023 7827 5049 7853
rect 7075 7827 7101 7853
rect 7127 7827 7153 7853
rect 7179 7827 7205 7853
rect 9231 7827 9257 7853
rect 9283 7827 9309 7853
rect 9335 7827 9361 7853
rect 1079 7743 1105 7769
rect 8359 7743 8385 7769
rect 1415 7687 1441 7713
rect 1471 7631 1497 7657
rect 2871 7631 2897 7657
rect 6399 7631 6425 7657
rect 6623 7631 6649 7657
rect 3207 7575 3233 7601
rect 4271 7575 4297 7601
rect 4943 7575 4969 7601
rect 6007 7575 6033 7601
rect 7015 7575 7041 7601
rect 8079 7575 8105 7601
rect 1685 7435 1711 7461
rect 1737 7435 1763 7461
rect 1789 7435 1815 7461
rect 3841 7435 3867 7461
rect 3893 7435 3919 7461
rect 3945 7435 3971 7461
rect 5997 7435 6023 7461
rect 6049 7435 6075 7461
rect 6101 7435 6127 7461
rect 8153 7435 8179 7461
rect 8205 7435 8231 7461
rect 8257 7435 8283 7461
rect 1415 7295 1441 7321
rect 3599 7295 3625 7321
rect 5559 7295 5585 7321
rect 7295 7295 7321 7321
rect 3151 7239 3177 7265
rect 3263 7239 3289 7265
rect 3431 7239 3457 7265
rect 3655 7239 3681 7265
rect 3767 7239 3793 7265
rect 4103 7239 4129 7265
rect 6063 7239 6089 7265
rect 6959 7239 6985 7265
rect 7071 7239 7097 7265
rect 7239 7239 7265 7265
rect 3039 7183 3065 7209
rect 4495 7183 4521 7209
rect 5727 7183 5753 7209
rect 5839 7183 5865 7209
rect 7351 7183 7377 7209
rect 7463 7183 7489 7209
rect 7575 7183 7601 7209
rect 7631 7183 7657 7209
rect 1471 7127 1497 7153
rect 3207 7127 3233 7153
rect 5895 7127 5921 7153
rect 2763 7043 2789 7069
rect 2815 7043 2841 7069
rect 2867 7043 2893 7069
rect 4919 7043 4945 7069
rect 4971 7043 4997 7069
rect 5023 7043 5049 7069
rect 7075 7043 7101 7069
rect 7127 7043 7153 7069
rect 7179 7043 7205 7069
rect 9231 7043 9257 7069
rect 9283 7043 9309 7069
rect 9335 7043 9361 7069
rect 3319 6959 3345 6985
rect 5111 6959 5137 6985
rect 5447 6959 5473 6985
rect 5727 6959 5753 6985
rect 5839 6959 5865 6985
rect 7071 6959 7097 6985
rect 1023 6903 1049 6929
rect 1471 6903 1497 6929
rect 2479 6903 2505 6929
rect 2647 6903 2673 6929
rect 2983 6903 3009 6929
rect 3655 6903 3681 6929
rect 3991 6903 4017 6929
rect 5223 6903 5249 6929
rect 5559 6903 5585 6929
rect 5615 6903 5641 6929
rect 6175 6903 6201 6929
rect 6959 6903 6985 6929
rect 855 6847 881 6873
rect 2871 6847 2897 6873
rect 3207 6847 3233 6873
rect 3543 6847 3569 6873
rect 3879 6847 3905 6873
rect 4999 6847 5025 6873
rect 5335 6847 5361 6873
rect 5895 6847 5921 6873
rect 6119 6847 6145 6873
rect 6511 6847 6537 6873
rect 6679 6847 6705 6873
rect 6903 6847 6929 6873
rect 1247 6791 1273 6817
rect 1415 6735 1441 6761
rect 1685 6651 1711 6677
rect 1737 6651 1763 6677
rect 1789 6651 1815 6677
rect 3841 6651 3867 6677
rect 3893 6651 3919 6677
rect 3945 6651 3971 6677
rect 5997 6651 6023 6677
rect 6049 6651 6075 6677
rect 6101 6651 6127 6677
rect 8153 6651 8179 6677
rect 8205 6651 8231 6677
rect 8257 6651 8283 6677
rect 5447 6567 5473 6593
rect 6791 6567 6817 6593
rect 2535 6511 2561 6537
rect 8975 6511 9001 6537
rect 1135 6455 1161 6481
rect 4551 6455 4577 6481
rect 5167 6455 5193 6481
rect 6735 6455 6761 6481
rect 7463 6455 7489 6481
rect 7575 6455 7601 6481
rect 8023 6455 8049 6481
rect 1471 6399 1497 6425
rect 5055 6399 5081 6425
rect 5615 6399 5641 6425
rect 5839 6399 5865 6425
rect 7239 6399 7265 6425
rect 7351 6399 7377 6425
rect 4663 6343 4689 6369
rect 6007 6343 6033 6369
rect 6847 6343 6873 6369
rect 6959 6343 6985 6369
rect 7463 6343 7489 6369
rect 2763 6259 2789 6285
rect 2815 6259 2841 6285
rect 2867 6259 2893 6285
rect 4919 6259 4945 6285
rect 4971 6259 4997 6285
rect 5023 6259 5049 6285
rect 7075 6259 7101 6285
rect 7127 6259 7153 6285
rect 7179 6259 7205 6285
rect 9231 6259 9257 6285
rect 9283 6259 9309 6285
rect 9335 6259 9361 6285
rect 1639 6175 1665 6201
rect 4495 6175 4521 6201
rect 4775 6175 4801 6201
rect 4831 6175 4857 6201
rect 6623 6175 6649 6201
rect 6903 6175 6929 6201
rect 7239 6175 7265 6201
rect 7687 6175 7713 6201
rect 7967 6175 7993 6201
rect 1303 6119 1329 6145
rect 1695 6119 1721 6145
rect 5223 6119 5249 6145
rect 6007 6119 6033 6145
rect 6119 6119 6145 6145
rect 6343 6119 6369 6145
rect 8023 6119 8049 6145
rect 1079 6063 1105 6089
rect 1415 6063 1441 6089
rect 1583 6063 1609 6089
rect 1975 6063 2001 6089
rect 2255 6063 2281 6089
rect 2367 6063 2393 6089
rect 3319 6063 3345 6089
rect 3487 6063 3513 6089
rect 4271 6063 4297 6089
rect 4383 6063 4409 6089
rect 4943 6063 4969 6089
rect 5111 6063 5137 6089
rect 5335 6063 5361 6089
rect 5615 6063 5641 6089
rect 5839 6063 5865 6089
rect 6063 6063 6089 6089
rect 6231 6063 6257 6089
rect 6847 6063 6873 6089
rect 7407 6063 7433 6089
rect 1359 6007 1385 6033
rect 3375 6007 3401 6033
rect 1191 5951 1217 5977
rect 1863 5951 1889 5977
rect 2199 5951 2225 5977
rect 4551 5951 4577 5977
rect 6511 5951 6537 5977
rect 6679 5951 6705 5977
rect 6903 5951 6929 5977
rect 7575 5951 7601 5977
rect 7743 5951 7769 5977
rect 7911 5951 7937 5977
rect 1685 5867 1711 5893
rect 1737 5867 1763 5893
rect 1789 5867 1815 5893
rect 3841 5867 3867 5893
rect 3893 5867 3919 5893
rect 3945 5867 3971 5893
rect 5997 5867 6023 5893
rect 6049 5867 6075 5893
rect 6101 5867 6127 5893
rect 8153 5867 8179 5893
rect 8205 5867 8231 5893
rect 8257 5867 8283 5893
rect 1471 5727 1497 5753
rect 2535 5727 2561 5753
rect 4103 5727 4129 5753
rect 6175 5727 6201 5753
rect 9087 5727 9113 5753
rect 1135 5671 1161 5697
rect 5839 5671 5865 5697
rect 6287 5671 6313 5697
rect 6847 5671 6873 5697
rect 7631 5671 7657 5697
rect 6735 5615 6761 5641
rect 6959 5615 6985 5641
rect 7127 5615 7153 5641
rect 8023 5615 8049 5641
rect 6455 5559 6481 5585
rect 7015 5559 7041 5585
rect 7183 5559 7209 5585
rect 7239 5559 7265 5585
rect 2763 5475 2789 5501
rect 2815 5475 2841 5501
rect 2867 5475 2893 5501
rect 4919 5475 4945 5501
rect 4971 5475 4997 5501
rect 5023 5475 5049 5501
rect 7075 5475 7101 5501
rect 7127 5475 7153 5501
rect 7179 5475 7205 5501
rect 9231 5475 9257 5501
rect 9283 5475 9309 5501
rect 9335 5475 9361 5501
rect 1247 5391 1273 5417
rect 4495 5391 4521 5417
rect 4887 5391 4913 5417
rect 8135 5391 8161 5417
rect 855 5335 881 5361
rect 1023 5335 1049 5361
rect 2199 5335 2225 5361
rect 2311 5335 2337 5361
rect 2647 5335 2673 5361
rect 4999 5335 5025 5361
rect 6175 5335 6201 5361
rect 2479 5279 2505 5305
rect 2815 5279 2841 5305
rect 4719 5279 4745 5305
rect 5167 5279 5193 5305
rect 7911 5279 7937 5305
rect 8079 5279 8105 5305
rect 8415 5279 8441 5305
rect 8695 5279 8721 5305
rect 1415 5223 1441 5249
rect 2143 5223 2169 5249
rect 3207 5223 3233 5249
rect 4271 5223 4297 5249
rect 4831 5223 4857 5249
rect 8303 5223 8329 5249
rect 8751 5223 8777 5249
rect 8975 5223 9001 5249
rect 1471 5167 1497 5193
rect 2479 5167 2505 5193
rect 8191 5167 8217 5193
rect 8919 5167 8945 5193
rect 1685 5083 1711 5109
rect 1737 5083 1763 5109
rect 1789 5083 1815 5109
rect 3841 5083 3867 5109
rect 3893 5083 3919 5109
rect 3945 5083 3971 5109
rect 5997 5083 6023 5109
rect 6049 5083 6075 5109
rect 6101 5083 6127 5109
rect 8153 5083 8179 5109
rect 8205 5083 8231 5109
rect 8257 5083 8283 5109
rect 3207 4999 3233 5025
rect 7127 4999 7153 5025
rect 2535 4943 2561 4969
rect 3543 4943 3569 4969
rect 4887 4943 4913 4969
rect 5615 4943 5641 4969
rect 6399 4943 6425 4969
rect 7239 4943 7265 4969
rect 7911 4943 7937 4969
rect 9031 4943 9057 4969
rect 1135 4887 1161 4913
rect 3263 4887 3289 4913
rect 4439 4887 4465 4913
rect 4831 4887 4857 4913
rect 5279 4887 5305 4913
rect 5447 4887 5473 4913
rect 6007 4887 6033 4913
rect 6287 4887 6313 4913
rect 6511 4887 6537 4913
rect 6903 4887 6929 4913
rect 7015 4887 7041 4913
rect 7351 4887 7377 4913
rect 7575 4887 7601 4913
rect 1471 4831 1497 4857
rect 2927 4831 2953 4857
rect 3039 4831 3065 4857
rect 4215 4831 4241 4857
rect 4775 4831 4801 4857
rect 5503 4831 5529 4857
rect 6175 4831 6201 4857
rect 3095 4775 3121 4801
rect 4047 4775 4073 4801
rect 4551 4775 4577 4801
rect 7407 4775 7433 4801
rect 2763 4691 2789 4717
rect 2815 4691 2841 4717
rect 2867 4691 2893 4717
rect 4919 4691 4945 4717
rect 4971 4691 4997 4717
rect 5023 4691 5049 4717
rect 7075 4691 7101 4717
rect 7127 4691 7153 4717
rect 7179 4691 7205 4717
rect 9231 4691 9257 4717
rect 9283 4691 9309 4717
rect 9335 4691 9361 4717
rect 1471 4607 1497 4633
rect 4383 4607 4409 4633
rect 4887 4607 4913 4633
rect 1023 4551 1049 4577
rect 1863 4551 1889 4577
rect 2031 4551 2057 4577
rect 2815 4551 2841 4577
rect 2983 4551 3009 4577
rect 3151 4551 3177 4577
rect 4495 4551 4521 4577
rect 5559 4551 5585 4577
rect 7575 4551 7601 4577
rect 8751 4551 8777 4577
rect 855 4495 881 4521
rect 1471 4495 1497 4521
rect 1695 4495 1721 4521
rect 2143 4495 2169 4521
rect 2367 4495 2393 4521
rect 3319 4495 3345 4521
rect 4271 4495 4297 4521
rect 4327 4495 4353 4521
rect 4831 4495 4857 4521
rect 4943 4495 4969 4521
rect 5111 4495 5137 4521
rect 5223 4495 5249 4521
rect 5447 4495 5473 4521
rect 6231 4495 6257 4521
rect 8695 4495 8721 4521
rect 8863 4495 8889 4521
rect 1247 4439 1273 4465
rect 2087 4439 2113 4465
rect 3207 4439 3233 4465
rect 5335 4439 5361 4465
rect 1639 4383 1665 4409
rect 2311 4383 2337 4409
rect 1685 4299 1711 4325
rect 1737 4299 1763 4325
rect 1789 4299 1815 4325
rect 3841 4299 3867 4325
rect 3893 4299 3919 4325
rect 3945 4299 3971 4325
rect 5997 4299 6023 4325
rect 6049 4299 6075 4325
rect 6101 4299 6127 4325
rect 8153 4299 8179 4325
rect 8205 4299 8231 4325
rect 8257 4299 8283 4325
rect 5447 4215 5473 4241
rect 6903 4215 6929 4241
rect 1471 4159 1497 4185
rect 2535 4159 2561 4185
rect 3823 4159 3849 4185
rect 4887 4159 4913 4185
rect 5055 4159 5081 4185
rect 6791 4159 6817 4185
rect 7855 4159 7881 4185
rect 8919 4159 8945 4185
rect 1135 4103 1161 4129
rect 3431 4103 3457 4129
rect 5335 4103 5361 4129
rect 5559 4103 5585 4129
rect 5783 4103 5809 4129
rect 6231 4103 6257 4129
rect 6343 4103 6369 4129
rect 6455 4103 6481 4129
rect 7519 4103 7545 4129
rect 5671 4047 5697 4073
rect 5895 4047 5921 4073
rect 5951 4047 5977 4073
rect 7071 4047 7097 4073
rect 6175 3991 6201 4017
rect 6287 3991 6313 4017
rect 6791 3991 6817 4017
rect 7239 3991 7265 4017
rect 2763 3907 2789 3933
rect 2815 3907 2841 3933
rect 2867 3907 2893 3933
rect 4919 3907 4945 3933
rect 4971 3907 4997 3933
rect 5023 3907 5049 3933
rect 7075 3907 7101 3933
rect 7127 3907 7153 3933
rect 7179 3907 7205 3933
rect 9231 3907 9257 3933
rect 9283 3907 9309 3933
rect 9335 3907 9361 3933
rect 1471 3823 1497 3849
rect 2703 3823 2729 3849
rect 3375 3823 3401 3849
rect 4495 3823 4521 3849
rect 5111 3823 5137 3849
rect 1415 3767 1441 3793
rect 3767 3767 3793 3793
rect 4719 3767 4745 3793
rect 4831 3767 4857 3793
rect 5335 3767 5361 3793
rect 6623 3767 6649 3793
rect 8863 3767 8889 3793
rect 2927 3711 2953 3737
rect 2983 3711 3009 3737
rect 3207 3711 3233 3737
rect 3319 3711 3345 3737
rect 3879 3711 3905 3737
rect 4215 3711 4241 3737
rect 4887 3711 4913 3737
rect 5055 3711 5081 3737
rect 6959 3711 6985 3737
rect 7351 3711 7377 3737
rect 8639 3711 8665 3737
rect 8975 3711 9001 3737
rect 2423 3655 2449 3681
rect 3095 3655 3121 3681
rect 8303 3655 8329 3681
rect 8751 3655 8777 3681
rect 1685 3515 1711 3541
rect 1737 3515 1763 3541
rect 1789 3515 1815 3541
rect 3841 3515 3867 3541
rect 3893 3515 3919 3541
rect 3945 3515 3971 3541
rect 5997 3515 6023 3541
rect 6049 3515 6075 3541
rect 6101 3515 6127 3541
rect 8153 3515 8179 3541
rect 8205 3515 8231 3541
rect 8257 3515 8283 3541
rect 4943 3431 4969 3457
rect 6231 3431 6257 3457
rect 3207 3375 3233 3401
rect 4271 3375 4297 3401
rect 5839 3375 5865 3401
rect 6791 3375 6817 3401
rect 8975 3375 9001 3401
rect 1415 3319 1441 3345
rect 1471 3319 1497 3345
rect 2871 3319 2897 3345
rect 4551 3319 4577 3345
rect 4999 3319 5025 3345
rect 5223 3319 5249 3345
rect 5783 3319 5809 3345
rect 6175 3319 6201 3345
rect 6399 3319 6425 3345
rect 7183 3319 7209 3345
rect 7519 3319 7545 3345
rect 7911 3319 7937 3345
rect 855 3263 881 3289
rect 1023 3263 1049 3289
rect 6735 3263 6761 3289
rect 6847 3263 6873 3289
rect 7071 3263 7097 3289
rect 1247 3207 1273 3233
rect 2763 3123 2789 3149
rect 2815 3123 2841 3149
rect 2867 3123 2893 3149
rect 4919 3123 4945 3149
rect 4971 3123 4997 3149
rect 5023 3123 5049 3149
rect 7075 3123 7101 3149
rect 7127 3123 7153 3149
rect 7179 3123 7205 3149
rect 9231 3123 9257 3149
rect 9283 3123 9309 3149
rect 9335 3123 9361 3149
rect 7183 3039 7209 3065
rect 7463 3039 7489 3065
rect 7743 3039 7769 3065
rect 8751 3039 8777 3065
rect 6511 2983 6537 3009
rect 8135 2983 8161 3009
rect 6903 2927 6929 2953
rect 7743 2927 7769 2953
rect 8191 2927 8217 2953
rect 5447 2871 5473 2897
rect 7071 2871 7097 2897
rect 7183 2871 7209 2897
rect 7407 2871 7433 2897
rect 1685 2731 1711 2757
rect 1737 2731 1763 2757
rect 1789 2731 1815 2757
rect 3841 2731 3867 2757
rect 3893 2731 3919 2757
rect 3945 2731 3971 2757
rect 5997 2731 6023 2757
rect 6049 2731 6075 2757
rect 6101 2731 6127 2757
rect 8153 2731 8179 2757
rect 8205 2731 8231 2757
rect 8257 2731 8283 2757
rect 2983 2647 3009 2673
rect 7295 2647 7321 2673
rect 6847 2591 6873 2617
rect 2927 2535 2953 2561
rect 7351 2535 7377 2561
rect 2763 2339 2789 2365
rect 2815 2339 2841 2365
rect 2867 2339 2893 2365
rect 4919 2339 4945 2365
rect 4971 2339 4997 2365
rect 5023 2339 5049 2365
rect 7075 2339 7101 2365
rect 7127 2339 7153 2365
rect 7179 2339 7205 2365
rect 9231 2339 9257 2365
rect 9283 2339 9309 2365
rect 9335 2339 9361 2365
rect 1023 2255 1049 2281
rect 855 2143 881 2169
rect 1247 2087 1273 2113
rect 1685 1947 1711 1973
rect 1737 1947 1763 1973
rect 1789 1947 1815 1973
rect 3841 1947 3867 1973
rect 3893 1947 3919 1973
rect 3945 1947 3971 1973
rect 5997 1947 6023 1973
rect 6049 1947 6075 1973
rect 6101 1947 6127 1973
rect 8153 1947 8179 1973
rect 8205 1947 8231 1973
rect 8257 1947 8283 1973
rect 967 1807 993 1833
rect 2143 1751 2169 1777
rect 8807 1695 8833 1721
rect 8919 1695 8945 1721
rect 9087 1695 9113 1721
rect 2763 1555 2789 1581
rect 2815 1555 2841 1581
rect 2867 1555 2893 1581
rect 4919 1555 4945 1581
rect 4971 1555 4997 1581
rect 5023 1555 5049 1581
rect 7075 1555 7101 1581
rect 7127 1555 7153 1581
rect 7179 1555 7205 1581
rect 9231 1555 9257 1581
rect 9283 1555 9309 1581
rect 9335 1555 9361 1581
<< metal2 >>
rect 2464 9600 2520 10000
rect 7392 9600 7448 10000
rect 1190 9226 1218 9231
rect 1190 8049 1218 9198
rect 1684 8246 1816 8251
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1684 8213 1816 8218
rect 1190 8023 1191 8049
rect 1217 8023 1218 8049
rect 854 7994 882 7999
rect 854 7947 882 7966
rect 1022 7938 1050 7943
rect 1022 7937 1162 7938
rect 1022 7911 1023 7937
rect 1049 7911 1162 7937
rect 1022 7910 1162 7911
rect 1022 7905 1050 7910
rect 1078 7770 1106 7775
rect 1078 7723 1106 7742
rect 1134 7546 1162 7910
rect 1190 7770 1218 8023
rect 1582 7994 1610 7999
rect 1582 7947 1610 7966
rect 1358 7938 1386 7943
rect 1358 7937 1442 7938
rect 1358 7911 1359 7937
rect 1385 7911 1442 7937
rect 1358 7910 1442 7911
rect 1358 7905 1386 7910
rect 1190 7737 1218 7742
rect 1414 7713 1442 7910
rect 1414 7687 1415 7713
rect 1441 7687 1442 7713
rect 1414 7681 1442 7687
rect 1470 7658 1498 7663
rect 1470 7611 1498 7630
rect 2478 7546 2506 9600
rect 3840 8246 3972 8251
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3840 8213 3972 8218
rect 5996 8246 6128 8251
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 5996 8213 6128 8218
rect 7406 8050 7434 9600
rect 7462 8666 7490 8671
rect 7462 8161 7490 8638
rect 8152 8246 8284 8251
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8152 8213 8284 8218
rect 7462 8135 7463 8161
rect 7489 8135 7490 8161
rect 7462 8129 7490 8135
rect 7406 8017 7434 8022
rect 8078 8049 8106 8055
rect 8078 8023 8079 8049
rect 8105 8023 8106 8049
rect 2762 7854 2894 7859
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2762 7821 2894 7826
rect 4918 7854 5050 7859
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 4918 7821 5050 7826
rect 7074 7854 7206 7859
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7074 7821 7206 7826
rect 2870 7657 2898 7663
rect 2870 7631 2871 7657
rect 2897 7631 2898 7657
rect 2870 7602 2898 7631
rect 2870 7569 2898 7574
rect 3150 7658 3178 7663
rect 1134 7518 1442 7546
rect 1414 7321 1442 7518
rect 2478 7513 2506 7518
rect 1684 7462 1816 7467
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1684 7429 1816 7434
rect 2982 7322 3010 7327
rect 1414 7295 1415 7321
rect 1441 7295 1442 7321
rect 1414 7289 1442 7295
rect 2926 7294 2982 7322
rect 1470 7154 1498 7159
rect 1470 7153 1610 7154
rect 1470 7127 1471 7153
rect 1497 7127 1610 7153
rect 1470 7126 1610 7127
rect 1470 7121 1498 7126
rect 1022 6930 1050 6935
rect 1470 6930 1498 6935
rect 1022 6929 1498 6930
rect 1022 6903 1023 6929
rect 1049 6903 1471 6929
rect 1497 6903 1498 6929
rect 1022 6902 1498 6903
rect 1022 6897 1050 6902
rect 1470 6897 1498 6902
rect 854 6873 882 6879
rect 854 6847 855 6873
rect 881 6847 882 6873
rect 854 6762 882 6847
rect 854 6729 882 6734
rect 1246 6817 1274 6823
rect 1246 6791 1247 6817
rect 1273 6791 1274 6817
rect 1246 6762 1274 6791
rect 1414 6762 1442 6767
rect 1246 6729 1274 6734
rect 1302 6761 1442 6762
rect 1302 6735 1415 6761
rect 1441 6735 1442 6761
rect 1302 6734 1442 6735
rect 1134 6481 1162 6487
rect 1134 6455 1135 6481
rect 1161 6455 1162 6481
rect 1078 6202 1106 6207
rect 1078 6089 1106 6174
rect 1078 6063 1079 6089
rect 1105 6063 1106 6089
rect 1078 6057 1106 6063
rect 1134 5697 1162 6455
rect 1302 6145 1330 6734
rect 1414 6729 1442 6734
rect 1582 6594 1610 7126
rect 2762 7070 2894 7075
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2762 7037 2894 7042
rect 2646 6986 2674 6991
rect 2478 6929 2506 6935
rect 2478 6903 2479 6929
rect 2505 6903 2506 6929
rect 1684 6678 1816 6683
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1684 6645 1816 6650
rect 1582 6566 1722 6594
rect 1470 6425 1498 6431
rect 1470 6399 1471 6425
rect 1497 6399 1498 6425
rect 1470 6202 1498 6399
rect 1638 6202 1666 6207
rect 1470 6201 1666 6202
rect 1470 6175 1639 6201
rect 1665 6175 1666 6201
rect 1470 6174 1666 6175
rect 1638 6169 1666 6174
rect 1302 6119 1303 6145
rect 1329 6119 1330 6145
rect 1302 6113 1330 6119
rect 1694 6145 1722 6566
rect 1694 6119 1695 6145
rect 1721 6119 1722 6145
rect 1694 6113 1722 6119
rect 1974 6202 2002 6207
rect 2478 6202 2506 6903
rect 2646 6929 2674 6958
rect 2646 6903 2647 6929
rect 2673 6903 2674 6929
rect 2646 6897 2674 6903
rect 2870 6874 2898 6879
rect 2926 6874 2954 7294
rect 2982 7289 3010 7294
rect 3150 7265 3178 7630
rect 6398 7658 6426 7663
rect 6622 7658 6650 7663
rect 6398 7657 6650 7658
rect 6398 7631 6399 7657
rect 6425 7631 6623 7657
rect 6649 7631 6650 7657
rect 6398 7630 6650 7631
rect 6398 7625 6426 7630
rect 3150 7239 3151 7265
rect 3177 7239 3178 7265
rect 3150 7233 3178 7239
rect 3206 7601 3234 7607
rect 3206 7575 3207 7601
rect 3233 7575 3234 7601
rect 3038 7210 3066 7215
rect 2702 6873 2954 6874
rect 2702 6847 2871 6873
rect 2897 6847 2954 6873
rect 2702 6846 2954 6847
rect 2982 7209 3066 7210
rect 2982 7183 3039 7209
rect 3065 7183 3066 7209
rect 2982 7182 3066 7183
rect 2982 6929 3010 7182
rect 3038 7177 3066 7182
rect 3206 7153 3234 7575
rect 4102 7602 4130 7607
rect 3840 7462 3972 7467
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3840 7429 3972 7434
rect 3598 7322 3626 7327
rect 3598 7275 3626 7294
rect 3766 7322 3794 7327
rect 3262 7266 3290 7271
rect 3262 7219 3290 7238
rect 3430 7265 3458 7271
rect 3430 7239 3431 7265
rect 3457 7239 3458 7265
rect 3206 7127 3207 7153
rect 3233 7127 3234 7153
rect 3206 7121 3234 7127
rect 3318 7210 3346 7215
rect 2982 6903 2983 6929
rect 3009 6903 3010 6929
rect 1414 6090 1442 6095
rect 1582 6090 1610 6095
rect 1414 6089 1582 6090
rect 1414 6063 1415 6089
rect 1441 6063 1582 6089
rect 1414 6062 1582 6063
rect 1414 6057 1442 6062
rect 1582 6043 1610 6062
rect 1974 6089 2002 6174
rect 2422 6174 2478 6202
rect 2254 6090 2282 6095
rect 1974 6063 1975 6089
rect 2001 6063 2002 6089
rect 1974 6057 2002 6063
rect 2142 6089 2282 6090
rect 2142 6063 2255 6089
rect 2281 6063 2282 6089
rect 2142 6062 2282 6063
rect 1358 6033 1386 6039
rect 1358 6007 1359 6033
rect 1385 6007 1386 6033
rect 1134 5671 1135 5697
rect 1161 5671 1162 5697
rect 854 5530 882 5535
rect 854 5361 882 5502
rect 1134 5418 1162 5671
rect 1190 5977 1218 5983
rect 1190 5951 1191 5977
rect 1217 5951 1218 5977
rect 1190 5586 1218 5951
rect 1358 5754 1386 6007
rect 1862 5978 1890 5983
rect 2142 5978 2170 6062
rect 2254 6057 2282 6062
rect 2366 6089 2394 6095
rect 2366 6063 2367 6089
rect 2393 6063 2394 6089
rect 1862 5977 2170 5978
rect 1862 5951 1863 5977
rect 1889 5951 2170 5977
rect 1862 5950 2170 5951
rect 2198 5978 2226 5983
rect 2198 5977 2338 5978
rect 2198 5951 2199 5977
rect 2225 5951 2338 5977
rect 2198 5950 2338 5951
rect 1862 5945 1890 5950
rect 2198 5945 2226 5950
rect 1684 5894 1816 5899
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1684 5861 1816 5866
rect 1470 5754 1498 5759
rect 1358 5753 1498 5754
rect 1358 5727 1471 5753
rect 1497 5727 1498 5753
rect 1358 5726 1498 5727
rect 1470 5721 1498 5726
rect 1190 5553 1218 5558
rect 2142 5586 2170 5591
rect 854 5335 855 5361
rect 881 5335 882 5361
rect 854 5329 882 5335
rect 1022 5361 1050 5367
rect 1022 5335 1023 5361
rect 1049 5335 1050 5361
rect 1022 5250 1050 5335
rect 1022 5217 1050 5222
rect 1134 4913 1162 5390
rect 1246 5530 1274 5535
rect 1246 5417 1274 5502
rect 1246 5391 1247 5417
rect 1273 5391 1274 5417
rect 1246 5385 1274 5391
rect 1414 5250 1442 5255
rect 1414 5203 1442 5222
rect 2142 5249 2170 5558
rect 2142 5223 2143 5249
rect 2169 5223 2170 5249
rect 2142 5217 2170 5223
rect 2198 5361 2226 5367
rect 2198 5335 2199 5361
rect 2225 5335 2226 5361
rect 1470 5193 1498 5199
rect 1470 5167 1471 5193
rect 1497 5167 1498 5193
rect 1470 4970 1498 5167
rect 2198 5194 2226 5335
rect 2310 5362 2338 5950
rect 2366 5922 2394 6063
rect 2366 5889 2394 5894
rect 2310 5315 2338 5334
rect 2198 5161 2226 5166
rect 1684 5110 1816 5115
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1684 5077 1816 5082
rect 1470 4937 1498 4942
rect 1638 5026 1666 5031
rect 1134 4887 1135 4913
rect 1161 4887 1162 4913
rect 1022 4577 1050 4583
rect 1022 4551 1023 4577
rect 1049 4551 1050 4577
rect 854 4521 882 4527
rect 854 4495 855 4521
rect 881 4495 882 4521
rect 854 4298 882 4495
rect 854 4265 882 4270
rect 1022 4214 1050 4551
rect 1022 4186 1106 4214
rect 1078 4018 1106 4186
rect 1134 4129 1162 4887
rect 1470 4857 1498 4863
rect 1470 4831 1471 4857
rect 1497 4831 1498 4857
rect 1470 4633 1498 4831
rect 1470 4607 1471 4633
rect 1497 4607 1498 4633
rect 1470 4601 1498 4607
rect 1414 4578 1442 4583
rect 1414 4522 1442 4550
rect 1470 4522 1498 4527
rect 1414 4521 1498 4522
rect 1414 4495 1471 4521
rect 1497 4495 1498 4521
rect 1414 4494 1498 4495
rect 1470 4489 1498 4494
rect 1526 4522 1554 4527
rect 1246 4465 1274 4471
rect 1246 4439 1247 4465
rect 1273 4439 1274 4465
rect 1246 4298 1274 4439
rect 1246 4265 1274 4270
rect 1470 4410 1498 4415
rect 1470 4185 1498 4382
rect 1470 4159 1471 4185
rect 1497 4159 1498 4185
rect 1470 4153 1498 4159
rect 1134 4103 1135 4129
rect 1161 4103 1162 4129
rect 1134 4097 1162 4103
rect 1078 3990 1442 4018
rect 1414 3793 1442 3990
rect 1470 3850 1498 3855
rect 1526 3850 1554 4494
rect 1638 4409 1666 4998
rect 1694 4970 1722 4975
rect 2422 4970 2450 6174
rect 2478 6169 2506 6174
rect 2534 6537 2562 6543
rect 2534 6511 2535 6537
rect 2561 6511 2562 6537
rect 2534 5922 2562 6511
rect 2534 5889 2562 5894
rect 2534 5754 2562 5759
rect 2534 5753 2618 5754
rect 2534 5727 2535 5753
rect 2561 5727 2618 5753
rect 2534 5726 2618 5727
rect 2534 5721 2562 5726
rect 2478 5306 2506 5311
rect 2478 5305 2562 5306
rect 2478 5279 2479 5305
rect 2505 5279 2562 5305
rect 2478 5278 2562 5279
rect 2478 5273 2506 5278
rect 2478 5193 2506 5199
rect 2478 5167 2479 5193
rect 2505 5167 2506 5193
rect 2478 5082 2506 5167
rect 2478 5049 2506 5054
rect 1694 4521 1722 4942
rect 2366 4942 2450 4970
rect 2534 4969 2562 5278
rect 2590 5194 2618 5726
rect 2590 5161 2618 5166
rect 2646 5362 2674 5367
rect 2646 5082 2674 5334
rect 2646 5049 2674 5054
rect 2534 4943 2535 4969
rect 2561 4943 2562 4969
rect 2030 4858 2058 4863
rect 1862 4578 1890 4583
rect 2030 4578 2058 4830
rect 1862 4577 2058 4578
rect 1862 4551 1863 4577
rect 1889 4551 2031 4577
rect 2057 4551 2058 4577
rect 1862 4550 2058 4551
rect 1862 4545 1890 4550
rect 2030 4545 2058 4550
rect 2366 4578 2394 4942
rect 2534 4914 2562 4943
rect 2534 4881 2562 4886
rect 1694 4495 1695 4521
rect 1721 4495 1722 4521
rect 1694 4489 1722 4495
rect 2142 4522 2170 4527
rect 2142 4475 2170 4494
rect 2366 4521 2394 4550
rect 2366 4495 2367 4521
rect 2393 4495 2394 4521
rect 2366 4489 2394 4495
rect 2422 4858 2450 4863
rect 1638 4383 1639 4409
rect 1665 4383 1666 4409
rect 1638 4377 1666 4383
rect 2086 4465 2114 4471
rect 2086 4439 2087 4465
rect 2113 4439 2114 4465
rect 2086 4410 2114 4439
rect 2086 4377 2114 4382
rect 2310 4410 2338 4415
rect 2310 4363 2338 4382
rect 1684 4326 1816 4331
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1684 4293 1816 4298
rect 1470 3849 1554 3850
rect 1470 3823 1471 3849
rect 1497 3823 1554 3849
rect 1470 3822 1554 3823
rect 1470 3817 1498 3822
rect 1414 3767 1415 3793
rect 1441 3767 1442 3793
rect 1414 3761 1442 3767
rect 2422 3681 2450 4830
rect 2702 4634 2730 6846
rect 2870 6841 2898 6846
rect 2762 6286 2894 6291
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2762 6253 2894 6258
rect 2982 6090 3010 6903
rect 3206 6986 3234 6991
rect 3318 6986 3346 7182
rect 3430 7098 3458 7239
rect 3654 7266 3682 7271
rect 3654 7219 3682 7238
rect 3766 7265 3794 7294
rect 3766 7239 3767 7265
rect 3793 7239 3794 7265
rect 3766 7233 3794 7239
rect 4102 7265 4130 7574
rect 4270 7601 4298 7607
rect 4270 7575 4271 7601
rect 4297 7575 4298 7601
rect 4270 7322 4298 7575
rect 4942 7601 4970 7607
rect 6006 7602 6034 7607
rect 4942 7575 4943 7601
rect 4969 7575 4970 7601
rect 4270 7289 4298 7294
rect 4438 7546 4466 7551
rect 4102 7239 4103 7265
rect 4129 7239 4130 7265
rect 3430 7070 3682 7098
rect 3206 6873 3234 6958
rect 3206 6847 3207 6873
rect 3233 6847 3234 6873
rect 3206 6841 3234 6847
rect 3262 6985 3346 6986
rect 3262 6959 3319 6985
rect 3345 6959 3346 6985
rect 3262 6958 3346 6959
rect 2982 6057 3010 6062
rect 2762 5502 2894 5507
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2762 5469 2894 5474
rect 2814 5418 2842 5423
rect 2814 5305 2842 5390
rect 2814 5279 2815 5305
rect 2841 5279 2842 5305
rect 2814 5273 2842 5279
rect 3206 5250 3234 5255
rect 3094 5249 3234 5250
rect 3094 5223 3207 5249
rect 3233 5223 3234 5249
rect 3094 5222 3234 5223
rect 2926 4858 2954 4863
rect 2926 4811 2954 4830
rect 3038 4857 3066 4863
rect 3038 4831 3039 4857
rect 3065 4831 3066 4857
rect 2762 4718 2894 4723
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 3038 4690 3066 4831
rect 3094 4801 3122 5222
rect 3206 5217 3234 5222
rect 3206 5138 3234 5143
rect 3094 4775 3095 4801
rect 3121 4775 3122 4801
rect 3094 4769 3122 4775
rect 3150 5082 3178 5087
rect 2762 4685 2894 4690
rect 2926 4662 3066 4690
rect 2702 4606 2842 4634
rect 2534 4522 2562 4527
rect 2534 4185 2562 4494
rect 2534 4159 2535 4185
rect 2561 4159 2562 4185
rect 2534 4153 2562 4159
rect 2702 3850 2730 4606
rect 2814 4577 2842 4606
rect 2814 4551 2815 4577
rect 2841 4551 2842 4577
rect 2814 4545 2842 4551
rect 2926 4214 2954 4662
rect 2982 4577 3010 4583
rect 2982 4551 2983 4577
rect 3009 4551 3010 4577
rect 2982 4522 3010 4551
rect 3150 4577 3178 5054
rect 3206 5025 3234 5110
rect 3206 4999 3207 5025
rect 3233 4999 3234 5025
rect 3206 4993 3234 4999
rect 3262 4970 3290 6958
rect 3318 6953 3346 6958
rect 3542 6986 3570 6991
rect 3542 6873 3570 6958
rect 3542 6847 3543 6873
rect 3569 6847 3570 6873
rect 3542 6841 3570 6847
rect 3654 6929 3682 7070
rect 3654 6903 3655 6929
rect 3681 6903 3682 6929
rect 3654 6482 3682 6903
rect 3878 6986 3906 6991
rect 3878 6873 3906 6958
rect 3878 6847 3879 6873
rect 3905 6847 3906 6873
rect 3878 6841 3906 6847
rect 3990 6929 4018 6935
rect 3990 6903 3991 6929
rect 4017 6903 4018 6929
rect 3990 6818 4018 6903
rect 3990 6785 4018 6790
rect 3840 6678 3972 6683
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3840 6645 3972 6650
rect 3654 6449 3682 6454
rect 3486 6202 3514 6207
rect 3318 6090 3346 6095
rect 3318 6043 3346 6062
rect 3486 6089 3514 6174
rect 3486 6063 3487 6089
rect 3513 6063 3514 6089
rect 3486 6057 3514 6063
rect 3374 6033 3402 6039
rect 3374 6007 3375 6033
rect 3401 6007 3402 6033
rect 3262 4913 3290 4942
rect 3262 4887 3263 4913
rect 3289 4887 3290 4913
rect 3262 4881 3290 4887
rect 3318 5922 3346 5927
rect 3318 4634 3346 5894
rect 3374 5138 3402 6007
rect 3840 5894 3972 5899
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3840 5861 3972 5866
rect 4102 5753 4130 7239
rect 4102 5727 4103 5753
rect 4129 5727 4130 5753
rect 3374 5105 3402 5110
rect 3430 5418 3458 5423
rect 3318 4601 3346 4606
rect 3150 4551 3151 4577
rect 3177 4551 3178 4577
rect 3150 4522 3178 4551
rect 2982 4494 3178 4522
rect 3318 4522 3346 4527
rect 3318 4475 3346 4494
rect 3206 4465 3234 4471
rect 3206 4439 3207 4465
rect 3233 4439 3234 4465
rect 3206 4410 3234 4439
rect 3206 4377 3234 4382
rect 2926 4186 3066 4214
rect 2926 4018 2954 4023
rect 2762 3934 2894 3939
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2762 3901 2894 3906
rect 2702 3803 2730 3822
rect 2926 3737 2954 3990
rect 2926 3711 2927 3737
rect 2953 3711 2954 3737
rect 2926 3705 2954 3711
rect 2982 3738 3010 3743
rect 2422 3655 2423 3681
rect 2449 3655 2450 3681
rect 1684 3542 1816 3547
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1684 3509 1816 3514
rect 1414 3346 1442 3351
rect 1022 3345 1442 3346
rect 1022 3319 1415 3345
rect 1441 3319 1442 3345
rect 1022 3318 1442 3319
rect 854 3289 882 3295
rect 854 3263 855 3289
rect 881 3263 882 3289
rect 854 3066 882 3263
rect 1022 3289 1050 3318
rect 1414 3313 1442 3318
rect 1470 3346 1498 3351
rect 1470 3299 1498 3318
rect 1022 3263 1023 3289
rect 1049 3263 1050 3289
rect 1022 3257 1050 3263
rect 854 3033 882 3038
rect 1246 3233 1274 3239
rect 1246 3207 1247 3233
rect 1273 3207 1274 3233
rect 1246 3066 1274 3207
rect 1246 3033 1274 3038
rect 1684 2758 1816 2763
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1684 2725 1816 2730
rect 1022 2562 1050 2567
rect 1022 2281 1050 2534
rect 1022 2255 1023 2281
rect 1049 2255 1050 2281
rect 1022 2249 1050 2255
rect 854 2169 882 2175
rect 854 2143 855 2169
rect 881 2143 882 2169
rect 854 2114 882 2143
rect 854 1834 882 2086
rect 1246 2114 1274 2119
rect 1246 2067 1274 2086
rect 1684 1974 1816 1979
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1684 1941 1816 1946
rect 854 1801 882 1806
rect 966 1833 994 1839
rect 966 1807 967 1833
rect 993 1807 994 1833
rect 966 658 994 1807
rect 2142 1778 2170 1783
rect 2422 1778 2450 3655
rect 2870 3626 2898 3631
rect 2870 3345 2898 3598
rect 2870 3319 2871 3345
rect 2897 3319 2898 3345
rect 2870 3313 2898 3319
rect 2762 3150 2894 3155
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2762 3117 2894 3122
rect 2982 2673 3010 3710
rect 3038 3346 3066 4186
rect 3430 4129 3458 5390
rect 4102 5418 4130 5727
rect 4102 5385 4130 5390
rect 4158 6818 4186 6823
rect 3840 5110 3972 5115
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3840 5077 3972 5082
rect 3542 4970 3570 4975
rect 3542 4923 3570 4942
rect 4046 4802 4074 4807
rect 4046 4755 4074 4774
rect 3840 4326 3972 4331
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3840 4293 3972 4298
rect 3822 4242 3850 4247
rect 3822 4185 3850 4214
rect 3822 4159 3823 4185
rect 3849 4159 3850 4185
rect 3822 4153 3850 4159
rect 3430 4103 3431 4129
rect 3457 4103 3458 4129
rect 3374 3850 3402 3855
rect 3374 3803 3402 3822
rect 3206 3794 3234 3799
rect 3206 3737 3234 3766
rect 3206 3711 3207 3737
rect 3233 3711 3234 3737
rect 3206 3705 3234 3711
rect 3318 3738 3346 3743
rect 3318 3691 3346 3710
rect 3094 3681 3122 3687
rect 3094 3655 3095 3681
rect 3121 3655 3122 3681
rect 3094 3458 3122 3655
rect 3430 3626 3458 4103
rect 4158 4018 4186 6790
rect 4214 6202 4242 6207
rect 4214 5250 4242 6174
rect 4270 6090 4298 6095
rect 4382 6090 4410 6095
rect 4270 6089 4354 6090
rect 4270 6063 4271 6089
rect 4297 6063 4354 6089
rect 4270 6062 4354 6063
rect 4270 6057 4298 6062
rect 4270 5250 4298 5255
rect 4214 5249 4298 5250
rect 4214 5223 4271 5249
rect 4297 5223 4298 5249
rect 4214 5222 4298 5223
rect 4270 5217 4298 5222
rect 4326 4970 4354 6062
rect 4382 6043 4410 6062
rect 4438 5418 4466 7518
rect 4494 7210 4522 7215
rect 4494 7163 4522 7182
rect 4942 7154 4970 7575
rect 5894 7601 6034 7602
rect 5894 7575 6007 7601
rect 6033 7575 6034 7601
rect 5894 7574 6034 7575
rect 5558 7321 5586 7327
rect 5558 7295 5559 7321
rect 5585 7295 5586 7321
rect 4942 7121 4970 7126
rect 5110 7210 5138 7215
rect 4918 7070 5050 7075
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 4918 7037 5050 7042
rect 5110 6985 5138 7182
rect 5446 6986 5474 6991
rect 5110 6959 5111 6985
rect 5137 6959 5138 6985
rect 5110 6953 5138 6959
rect 5278 6985 5474 6986
rect 5278 6959 5447 6985
rect 5473 6959 5474 6985
rect 5278 6958 5474 6959
rect 5222 6930 5250 6935
rect 5278 6930 5306 6958
rect 5446 6953 5474 6958
rect 5222 6929 5306 6930
rect 5222 6903 5223 6929
rect 5249 6903 5306 6929
rect 5222 6902 5306 6903
rect 5558 6929 5586 7295
rect 5726 7210 5754 7215
rect 5838 7210 5866 7215
rect 5670 7209 5754 7210
rect 5670 7183 5727 7209
rect 5753 7183 5754 7209
rect 5670 7182 5754 7183
rect 5558 6903 5559 6929
rect 5585 6903 5586 6929
rect 5222 6897 5250 6902
rect 4998 6874 5026 6879
rect 4774 6873 5026 6874
rect 4774 6847 4999 6873
rect 5025 6847 5026 6873
rect 4774 6846 5026 6847
rect 4550 6481 4578 6487
rect 4550 6455 4551 6481
rect 4577 6455 4578 6481
rect 4494 6202 4522 6207
rect 4494 6155 4522 6174
rect 4550 6146 4578 6455
rect 4662 6370 4690 6375
rect 4662 6323 4690 6342
rect 4774 6201 4802 6846
rect 4998 6841 5026 6846
rect 5166 6874 5194 6879
rect 5166 6481 5194 6846
rect 5166 6455 5167 6481
rect 5193 6455 5194 6481
rect 5054 6426 5082 6431
rect 5054 6379 5082 6398
rect 4918 6286 5050 6291
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 4918 6253 5050 6258
rect 4774 6175 4775 6201
rect 4801 6175 4802 6201
rect 4774 6169 4802 6175
rect 4830 6202 4858 6207
rect 4830 6155 4858 6174
rect 4550 6113 4578 6118
rect 4886 6146 4914 6151
rect 4550 5977 4578 5983
rect 4550 5951 4551 5977
rect 4577 5951 4578 5977
rect 4550 5586 4578 5951
rect 4886 5586 4914 6118
rect 4942 6090 4970 6095
rect 4942 6043 4970 6062
rect 5110 6089 5138 6095
rect 5110 6063 5111 6089
rect 5137 6063 5138 6089
rect 5110 6034 5138 6063
rect 5110 6001 5138 6006
rect 4550 5553 4578 5558
rect 4830 5558 4914 5586
rect 4494 5418 4522 5423
rect 4438 5390 4494 5418
rect 4830 5418 4858 5558
rect 5166 5530 5194 6455
rect 5334 6873 5362 6879
rect 5334 6847 5335 6873
rect 5361 6847 5362 6873
rect 5334 6818 5362 6847
rect 5334 6426 5362 6790
rect 5446 6594 5474 6599
rect 5558 6594 5586 6903
rect 5614 6930 5642 6935
rect 5614 6883 5642 6902
rect 5446 6593 5586 6594
rect 5446 6567 5447 6593
rect 5473 6567 5586 6593
rect 5446 6566 5586 6567
rect 5446 6561 5474 6566
rect 5670 6538 5698 7182
rect 5726 7177 5754 7182
rect 5782 7209 5866 7210
rect 5782 7183 5839 7209
rect 5865 7183 5866 7209
rect 5782 7182 5866 7183
rect 5726 6986 5754 6991
rect 5782 6986 5810 7182
rect 5838 7177 5866 7182
rect 5894 7153 5922 7574
rect 6006 7569 6034 7574
rect 5996 7462 6128 7467
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 5996 7429 6128 7434
rect 6174 7322 6202 7327
rect 5894 7127 5895 7153
rect 5921 7127 5922 7153
rect 5894 7121 5922 7127
rect 6062 7265 6090 7271
rect 6062 7239 6063 7265
rect 6089 7239 6090 7265
rect 5726 6985 5810 6986
rect 5726 6959 5727 6985
rect 5753 6959 5810 6985
rect 5726 6958 5810 6959
rect 5838 7098 5866 7103
rect 5838 6985 5866 7070
rect 5838 6959 5839 6985
rect 5865 6959 5866 6985
rect 5726 6953 5754 6958
rect 5838 6953 5866 6959
rect 5894 6873 5922 6879
rect 5894 6847 5895 6873
rect 5921 6847 5922 6873
rect 5894 6762 5922 6847
rect 6062 6762 6090 7239
rect 6174 6929 6202 7294
rect 6174 6903 6175 6929
rect 6201 6903 6202 6929
rect 6174 6897 6202 6903
rect 6510 7098 6538 7103
rect 6118 6874 6146 6879
rect 6118 6827 6146 6846
rect 6510 6873 6538 7070
rect 6510 6847 6511 6873
rect 6537 6847 6538 6873
rect 6510 6841 6538 6847
rect 6062 6734 6202 6762
rect 5894 6729 5922 6734
rect 5996 6678 6128 6683
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 5996 6645 6128 6650
rect 6174 6594 6202 6734
rect 6174 6561 6202 6566
rect 5558 6510 5698 6538
rect 5558 6426 5586 6510
rect 5334 6398 5586 6426
rect 5222 6146 5250 6151
rect 5222 6099 5250 6118
rect 5334 6089 5362 6095
rect 5334 6063 5335 6089
rect 5361 6063 5362 6089
rect 5334 5922 5362 6063
rect 5334 5889 5362 5894
rect 4918 5502 5050 5507
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 4918 5469 5050 5474
rect 5110 5502 5194 5530
rect 5222 5586 5250 5591
rect 4886 5418 4914 5423
rect 4830 5417 4914 5418
rect 4830 5391 4887 5417
rect 4913 5391 4914 5417
rect 4830 5390 4914 5391
rect 4494 5371 4522 5390
rect 4718 5306 4746 5311
rect 4214 4858 4242 4863
rect 4326 4858 4354 4942
rect 4214 4857 4354 4858
rect 4214 4831 4215 4857
rect 4241 4831 4354 4857
rect 4214 4830 4354 4831
rect 4382 5305 4746 5306
rect 4382 5279 4719 5305
rect 4745 5279 4746 5305
rect 4382 5278 4746 5279
rect 4214 4825 4242 4830
rect 4382 4802 4410 5278
rect 4718 5273 4746 5278
rect 4830 5250 4858 5255
rect 4830 5203 4858 5222
rect 4718 5194 4746 5199
rect 4382 4633 4410 4774
rect 4438 4913 4466 4919
rect 4438 4887 4439 4913
rect 4465 4887 4466 4913
rect 4438 4746 4466 4887
rect 4438 4713 4466 4718
rect 4494 4802 4522 4807
rect 4382 4607 4383 4633
rect 4409 4607 4410 4633
rect 4382 4601 4410 4607
rect 4494 4577 4522 4774
rect 4494 4551 4495 4577
rect 4521 4551 4522 4577
rect 4270 4521 4298 4527
rect 4270 4495 4271 4521
rect 4297 4495 4298 4521
rect 4158 3985 4186 3990
rect 4214 4466 4242 4471
rect 3430 3593 3458 3598
rect 3766 3793 3794 3799
rect 3766 3767 3767 3793
rect 3793 3767 3794 3793
rect 3766 3626 3794 3767
rect 3878 3738 3906 3743
rect 3878 3691 3906 3710
rect 4214 3737 4242 4438
rect 4270 4186 4298 4495
rect 4326 4522 4354 4527
rect 4326 4475 4354 4494
rect 4494 4522 4522 4551
rect 4550 4801 4578 4807
rect 4550 4775 4551 4801
rect 4577 4775 4578 4801
rect 4550 4578 4578 4775
rect 4550 4545 4578 4550
rect 4494 4489 4522 4494
rect 4718 4410 4746 5166
rect 4886 4969 4914 5390
rect 4886 4943 4887 4969
rect 4913 4943 4914 4969
rect 4886 4937 4914 4943
rect 4998 5361 5026 5367
rect 4998 5335 4999 5361
rect 5025 5335 5026 5361
rect 4830 4914 4858 4919
rect 4830 4867 4858 4886
rect 4774 4858 4802 4863
rect 4774 4811 4802 4830
rect 4998 4802 5026 5335
rect 4830 4774 5026 4802
rect 4830 4746 4858 4774
rect 4830 4634 4858 4718
rect 4918 4718 5050 4723
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 4918 4685 5050 4690
rect 4886 4634 4914 4639
rect 5110 4634 5138 5502
rect 5166 5418 5194 5423
rect 5166 5305 5194 5390
rect 5166 5279 5167 5305
rect 5193 5279 5194 5305
rect 5166 5273 5194 5279
rect 4830 4633 4914 4634
rect 4830 4607 4887 4633
rect 4913 4607 4914 4633
rect 4830 4606 4914 4607
rect 4886 4601 4914 4606
rect 5054 4606 5138 4634
rect 4830 4522 4858 4527
rect 4830 4475 4858 4494
rect 4942 4521 4970 4527
rect 4942 4495 4943 4521
rect 4969 4495 4970 4521
rect 4942 4410 4970 4495
rect 4718 4382 4970 4410
rect 5054 4298 5082 4606
rect 4270 4153 4298 4158
rect 4886 4186 4914 4191
rect 4886 4139 4914 4158
rect 5054 4185 5082 4270
rect 5054 4159 5055 4185
rect 5081 4159 5082 4185
rect 5054 4153 5082 4159
rect 5110 4521 5138 4527
rect 5110 4495 5111 4521
rect 5137 4495 5138 4521
rect 5110 4130 5138 4495
rect 5222 4521 5250 5558
rect 5222 4495 5223 4521
rect 5249 4495 5250 4521
rect 5222 4489 5250 4495
rect 5278 4913 5306 4919
rect 5278 4887 5279 4913
rect 5305 4887 5306 4913
rect 5278 4858 5306 4887
rect 5446 4914 5474 4919
rect 5446 4867 5474 4886
rect 5278 4578 5306 4830
rect 5502 4857 5530 4863
rect 5502 4831 5503 4857
rect 5529 4831 5530 4857
rect 5502 4634 5530 4831
rect 5502 4601 5530 4606
rect 5278 4550 5418 4578
rect 5278 4298 5306 4550
rect 5110 4097 5138 4102
rect 5166 4270 5306 4298
rect 5334 4465 5362 4471
rect 5334 4439 5335 4465
rect 5361 4439 5362 4465
rect 4918 3934 5050 3939
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 4918 3901 5050 3906
rect 4494 3850 4522 3855
rect 5110 3850 5138 3855
rect 4522 3822 4578 3850
rect 4494 3803 4522 3822
rect 4214 3711 4215 3737
rect 4241 3711 4242 3737
rect 4214 3705 4242 3711
rect 3766 3593 3794 3598
rect 4270 3626 4298 3631
rect 3840 3542 3972 3547
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3840 3509 3972 3514
rect 3094 3430 3234 3458
rect 3206 3401 3234 3430
rect 3206 3375 3207 3401
rect 3233 3375 3234 3401
rect 3206 3369 3234 3375
rect 4270 3401 4298 3598
rect 4270 3375 4271 3401
rect 4297 3375 4298 3401
rect 4270 3369 4298 3375
rect 3038 3313 3066 3318
rect 4550 3345 4578 3822
rect 5110 3803 5138 3822
rect 4718 3794 4746 3799
rect 4718 3747 4746 3766
rect 4830 3793 4858 3799
rect 4830 3767 4831 3793
rect 4857 3767 4858 3793
rect 4830 3626 4858 3767
rect 4886 3738 4914 3743
rect 5054 3738 5082 3743
rect 5166 3738 5194 4270
rect 5334 4242 5362 4439
rect 5390 4242 5418 4550
rect 5558 4577 5586 6398
rect 5614 6426 5642 6431
rect 5614 6425 5698 6426
rect 5614 6399 5615 6425
rect 5641 6399 5698 6425
rect 5614 6398 5698 6399
rect 5614 6393 5642 6398
rect 5614 6202 5642 6207
rect 5614 6089 5642 6174
rect 5614 6063 5615 6089
rect 5641 6063 5642 6089
rect 5614 4969 5642 6063
rect 5670 6090 5698 6398
rect 5838 6425 5866 6431
rect 5838 6399 5839 6425
rect 5865 6399 5866 6425
rect 5838 6202 5866 6399
rect 6006 6369 6034 6375
rect 6006 6343 6007 6369
rect 6033 6343 6034 6369
rect 5838 6169 5866 6174
rect 5950 6314 5978 6319
rect 5838 6090 5866 6095
rect 5670 6089 5866 6090
rect 5670 6063 5839 6089
rect 5865 6063 5866 6089
rect 5670 6062 5866 6063
rect 5670 6034 5698 6062
rect 5838 6057 5866 6062
rect 5670 6001 5698 6006
rect 5950 5978 5978 6286
rect 6006 6258 6034 6343
rect 6342 6370 6370 6375
rect 6006 6230 6202 6258
rect 6006 6146 6034 6151
rect 6006 6099 6034 6118
rect 6118 6145 6146 6151
rect 6118 6119 6119 6145
rect 6145 6119 6146 6145
rect 6062 6090 6090 6095
rect 6062 6043 6090 6062
rect 6118 5978 6146 6119
rect 5894 5950 6146 5978
rect 6174 6090 6202 6230
rect 6342 6146 6370 6342
rect 6286 6145 6370 6146
rect 6286 6119 6343 6145
rect 6369 6119 6370 6145
rect 6286 6118 6370 6119
rect 6230 6090 6258 6095
rect 6174 6062 6230 6090
rect 5894 5922 5922 5950
rect 5838 5697 5866 5703
rect 5838 5671 5839 5697
rect 5865 5671 5866 5697
rect 5838 5362 5866 5671
rect 5838 5329 5866 5334
rect 5614 4943 5615 4969
rect 5641 4943 5642 4969
rect 5614 4937 5642 4943
rect 5558 4551 5559 4577
rect 5585 4551 5586 4577
rect 5558 4545 5586 4551
rect 5894 4578 5922 5894
rect 5996 5894 6128 5899
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 5996 5861 6128 5866
rect 6174 5753 6202 6062
rect 6230 6043 6258 6062
rect 6286 5810 6314 6118
rect 6342 6113 6370 6118
rect 6174 5727 6175 5753
rect 6201 5727 6202 5753
rect 6174 5721 6202 5727
rect 6230 5782 6314 5810
rect 6510 5977 6538 5983
rect 6510 5951 6511 5977
rect 6537 5951 6538 5977
rect 6230 5586 6258 5782
rect 6286 5698 6314 5703
rect 6286 5697 6370 5698
rect 6286 5671 6287 5697
rect 6313 5671 6370 5697
rect 6286 5670 6370 5671
rect 6286 5665 6314 5670
rect 6230 5558 6314 5586
rect 6174 5362 6202 5367
rect 6202 5334 6258 5362
rect 6174 5315 6202 5334
rect 5996 5110 6128 5115
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 5996 5077 6128 5082
rect 5894 4545 5922 4550
rect 6006 4913 6034 4919
rect 6006 4887 6007 4913
rect 6033 4887 6034 4913
rect 5446 4522 5474 4527
rect 5446 4521 5530 4522
rect 5446 4495 5447 4521
rect 5473 4495 5530 4521
rect 5446 4494 5530 4495
rect 5446 4489 5474 4494
rect 5502 4410 5530 4494
rect 6006 4410 6034 4887
rect 6174 4857 6202 4863
rect 6174 4831 6175 4857
rect 6201 4831 6202 4857
rect 6174 4578 6202 4831
rect 6174 4545 6202 4550
rect 6230 4521 6258 5334
rect 6286 4913 6314 5558
rect 6286 4887 6287 4913
rect 6313 4887 6314 4913
rect 6286 4881 6314 4887
rect 6342 5250 6370 5670
rect 6230 4495 6231 4521
rect 6257 4495 6258 4521
rect 6230 4489 6258 4495
rect 5502 4382 5810 4410
rect 5726 4298 5754 4303
rect 5446 4242 5474 4247
rect 5390 4241 5474 4242
rect 5390 4215 5447 4241
rect 5473 4215 5474 4241
rect 5390 4214 5474 4215
rect 5334 4209 5362 4214
rect 5446 4209 5474 4214
rect 5222 4186 5250 4191
rect 5670 4186 5698 4191
rect 5250 4158 5306 4186
rect 5222 4153 5250 4158
rect 5278 4130 5306 4158
rect 5334 4130 5362 4135
rect 5278 4129 5362 4130
rect 5278 4103 5335 4129
rect 5361 4103 5362 4129
rect 5278 4102 5362 4103
rect 5334 4074 5362 4102
rect 5334 3793 5362 4046
rect 5334 3767 5335 3793
rect 5361 3767 5362 3793
rect 5334 3761 5362 3767
rect 5558 4130 5586 4135
rect 5558 3794 5586 4102
rect 5670 4074 5698 4158
rect 5558 3761 5586 3766
rect 5614 4073 5698 4074
rect 5614 4047 5671 4073
rect 5697 4047 5698 4073
rect 5614 4046 5698 4047
rect 4914 3710 4970 3738
rect 4886 3691 4914 3710
rect 4830 3593 4858 3598
rect 4942 3457 4970 3710
rect 5054 3737 5194 3738
rect 5054 3711 5055 3737
rect 5081 3711 5194 3737
rect 5054 3710 5194 3711
rect 5054 3705 5082 3710
rect 4942 3431 4943 3457
rect 4969 3431 4970 3457
rect 4942 3425 4970 3431
rect 4550 3319 4551 3345
rect 4577 3319 4578 3345
rect 4550 3313 4578 3319
rect 4998 3346 5026 3351
rect 4998 3299 5026 3318
rect 5222 3345 5250 3351
rect 5222 3319 5223 3345
rect 5249 3319 5250 3345
rect 5222 3290 5250 3319
rect 5222 3257 5250 3262
rect 4918 3150 5050 3155
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 4918 3117 5050 3122
rect 5446 2898 5474 2903
rect 5614 2898 5642 4046
rect 5670 4041 5698 4046
rect 5726 3962 5754 4270
rect 5782 4129 5810 4382
rect 5894 4382 6034 4410
rect 5894 4186 5922 4382
rect 5996 4326 6128 4331
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 5996 4293 6128 4298
rect 6342 4214 6370 5222
rect 6398 5642 6426 5647
rect 6398 4969 6426 5614
rect 6454 5585 6482 5591
rect 6454 5559 6455 5585
rect 6481 5559 6482 5585
rect 6454 5026 6482 5559
rect 6454 4993 6482 4998
rect 6398 4943 6399 4969
rect 6425 4943 6426 4969
rect 6398 4937 6426 4943
rect 6510 4970 6538 5951
rect 6566 5754 6594 7630
rect 6622 7625 6650 7630
rect 7014 7602 7042 7607
rect 8078 7602 8106 8023
rect 8358 8050 8386 8055
rect 8358 7769 8386 8022
rect 8582 8050 8610 8055
rect 8582 8003 8610 8022
rect 8358 7743 8359 7769
rect 8385 7743 8386 7769
rect 8358 7737 8386 7743
rect 8470 7937 8498 7943
rect 8470 7911 8471 7937
rect 8497 7911 8498 7937
rect 7014 7601 7322 7602
rect 7014 7575 7015 7601
rect 7041 7575 7322 7601
rect 7014 7574 7322 7575
rect 7014 7569 7042 7574
rect 7294 7321 7322 7574
rect 7294 7295 7295 7321
rect 7321 7295 7322 7321
rect 7294 7289 7322 7295
rect 7574 7601 8106 7602
rect 7574 7575 8079 7601
rect 8105 7575 8106 7601
rect 7574 7574 8106 7575
rect 6958 7266 6986 7271
rect 7070 7266 7098 7271
rect 6986 7265 7098 7266
rect 6986 7239 7071 7265
rect 7097 7239 7098 7265
rect 6986 7238 7098 7239
rect 6958 7219 6986 7238
rect 7070 7233 7098 7238
rect 7238 7265 7266 7271
rect 7238 7239 7239 7265
rect 7265 7239 7266 7265
rect 7074 7070 7206 7075
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7074 7037 7206 7042
rect 7070 6986 7098 6991
rect 7238 6986 7266 7239
rect 7518 7266 7546 7271
rect 7350 7210 7378 7215
rect 7462 7210 7490 7215
rect 7350 7209 7490 7210
rect 7350 7183 7351 7209
rect 7377 7183 7463 7209
rect 7489 7183 7490 7209
rect 7350 7182 7490 7183
rect 7350 7177 7378 7182
rect 7462 7177 7490 7182
rect 7070 6985 7266 6986
rect 7070 6959 7071 6985
rect 7097 6959 7266 6985
rect 7070 6958 7266 6959
rect 7070 6953 7098 6958
rect 6958 6930 6986 6935
rect 6958 6929 7042 6930
rect 6958 6903 6959 6929
rect 6985 6903 7042 6929
rect 6958 6902 7042 6903
rect 6958 6897 6986 6902
rect 6678 6874 6706 6879
rect 6902 6874 6930 6879
rect 6678 6873 6930 6874
rect 6678 6847 6679 6873
rect 6705 6847 6903 6873
rect 6929 6847 6930 6873
rect 6678 6846 6930 6847
rect 6678 6841 6706 6846
rect 6734 6481 6762 6846
rect 6902 6841 6930 6846
rect 6790 6594 6818 6599
rect 6790 6547 6818 6566
rect 6734 6455 6735 6481
rect 6761 6455 6762 6481
rect 6734 6449 6762 6455
rect 6566 5721 6594 5726
rect 6622 6370 6650 6375
rect 6846 6370 6874 6375
rect 6622 6201 6650 6342
rect 6622 6175 6623 6201
rect 6649 6175 6650 6201
rect 6622 5698 6650 6175
rect 6790 6342 6846 6370
rect 6734 6146 6762 6151
rect 6790 6146 6818 6342
rect 6846 6323 6874 6342
rect 6958 6369 6986 6375
rect 6958 6343 6959 6369
rect 6985 6343 6986 6369
rect 6902 6314 6930 6319
rect 6902 6201 6930 6286
rect 6902 6175 6903 6201
rect 6929 6175 6930 6201
rect 6902 6169 6930 6175
rect 6762 6118 6818 6146
rect 6734 6113 6762 6118
rect 6846 6090 6874 6095
rect 6678 5978 6706 5983
rect 6678 5931 6706 5950
rect 6846 5922 6874 6062
rect 6958 6090 6986 6343
rect 7014 6202 7042 6902
rect 7462 6482 7490 6487
rect 7462 6435 7490 6454
rect 7238 6425 7266 6431
rect 7238 6399 7239 6425
rect 7265 6399 7266 6425
rect 7238 6370 7266 6399
rect 7238 6337 7266 6342
rect 7350 6425 7378 6431
rect 7350 6399 7351 6425
rect 7377 6399 7378 6425
rect 7074 6286 7206 6291
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7074 6253 7206 6258
rect 7014 6169 7042 6174
rect 7238 6202 7266 6207
rect 7350 6202 7378 6399
rect 7266 6174 7378 6202
rect 7462 6369 7490 6375
rect 7462 6343 7463 6369
rect 7489 6343 7490 6369
rect 7238 6155 7266 6174
rect 6958 6057 6986 6062
rect 7406 6090 7434 6095
rect 7406 6043 7434 6062
rect 6734 5894 6874 5922
rect 6902 5977 6930 5983
rect 6902 5951 6903 5977
rect 6929 5951 6930 5977
rect 6734 5866 6762 5894
rect 6622 5665 6650 5670
rect 6678 5838 6762 5866
rect 6510 4913 6538 4942
rect 6510 4887 6511 4913
rect 6537 4887 6538 4913
rect 6510 4881 6538 4887
rect 6678 4802 6706 5838
rect 6790 5810 6818 5815
rect 6734 5641 6762 5647
rect 6734 5615 6735 5641
rect 6761 5615 6762 5641
rect 6734 4970 6762 5615
rect 6734 4937 6762 4942
rect 6790 4858 6818 5782
rect 6846 5698 6874 5703
rect 6846 5651 6874 5670
rect 6902 5642 6930 5951
rect 6958 5642 6986 5647
rect 6902 5641 6986 5642
rect 6902 5615 6959 5641
rect 6985 5615 6986 5641
rect 6902 5614 6986 5615
rect 6958 5609 6986 5614
rect 7126 5642 7154 5647
rect 7126 5595 7154 5614
rect 7462 5642 7490 6343
rect 7462 5609 7490 5614
rect 7014 5585 7042 5591
rect 7014 5559 7015 5585
rect 7041 5559 7042 5585
rect 6958 5530 6986 5535
rect 6902 5502 6958 5530
rect 6902 4913 6930 5502
rect 6958 5497 6986 5502
rect 7014 5306 7042 5559
rect 7182 5586 7210 5605
rect 7182 5553 7210 5558
rect 7238 5586 7266 5591
rect 7238 5585 7322 5586
rect 7238 5559 7239 5585
rect 7265 5559 7322 5585
rect 7238 5558 7322 5559
rect 7238 5553 7266 5558
rect 7074 5502 7206 5507
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7074 5469 7206 5474
rect 7014 5273 7042 5278
rect 6902 4887 6903 4913
rect 6929 4887 6930 4913
rect 6902 4881 6930 4887
rect 7014 5026 7042 5031
rect 7014 4913 7042 4998
rect 7126 5026 7154 5031
rect 7126 4979 7154 4998
rect 7014 4887 7015 4913
rect 7041 4887 7042 4913
rect 7014 4881 7042 4887
rect 7238 4970 7266 4975
rect 6678 4769 6706 4774
rect 6734 4830 6818 4858
rect 5894 4153 5922 4158
rect 6286 4186 6370 4214
rect 6622 4186 6650 4191
rect 5782 4103 5783 4129
rect 5809 4103 5810 4129
rect 5782 4097 5810 4103
rect 6230 4130 6258 4135
rect 6286 4130 6314 4186
rect 6342 4130 6370 4135
rect 6286 4129 6370 4130
rect 6286 4103 6343 4129
rect 6369 4103 6370 4129
rect 6286 4102 6370 4103
rect 6230 4083 6258 4102
rect 6342 4097 6370 4102
rect 6454 4130 6482 4135
rect 6454 4083 6482 4102
rect 5894 4074 5922 4079
rect 5894 4027 5922 4046
rect 5950 4073 5978 4079
rect 5950 4047 5951 4073
rect 5977 4047 5978 4073
rect 5950 4018 5978 4047
rect 6174 4018 6202 4023
rect 5950 4017 6202 4018
rect 5950 3991 6175 4017
rect 6201 3991 6202 4017
rect 5950 3990 6202 3991
rect 5726 3934 5810 3962
rect 5446 2897 5642 2898
rect 5446 2871 5447 2897
rect 5473 2871 5642 2897
rect 5446 2870 5642 2871
rect 5782 3345 5810 3934
rect 6174 3850 6202 3990
rect 6174 3817 6202 3822
rect 6286 4017 6314 4023
rect 6286 3991 6287 4017
rect 6313 3991 6314 4017
rect 5838 3626 5866 3631
rect 5838 3401 5866 3598
rect 5996 3542 6128 3547
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 5996 3509 6128 3514
rect 6230 3458 6258 3463
rect 6230 3411 6258 3430
rect 5838 3375 5839 3401
rect 5865 3375 5866 3401
rect 5838 3369 5866 3375
rect 6286 3402 6314 3991
rect 6622 3793 6650 4158
rect 6734 3850 6762 4830
rect 6902 4802 6930 4807
rect 6846 4634 6874 4639
rect 6790 4185 6818 4191
rect 6790 4159 6791 4185
rect 6817 4159 6818 4185
rect 6790 4130 6818 4159
rect 6790 4097 6818 4102
rect 6790 4017 6818 4023
rect 6790 3991 6791 4017
rect 6817 3991 6818 4017
rect 6790 3962 6818 3991
rect 6790 3929 6818 3934
rect 6734 3817 6762 3822
rect 6622 3767 6623 3793
rect 6649 3767 6650 3793
rect 6622 3761 6650 3767
rect 6790 3402 6818 3407
rect 6286 3369 6314 3374
rect 6510 3401 6818 3402
rect 6510 3375 6791 3401
rect 6817 3375 6818 3401
rect 6510 3374 6818 3375
rect 5782 3319 5783 3345
rect 5809 3319 5810 3345
rect 5782 2898 5810 3319
rect 5446 2865 5474 2870
rect 5782 2865 5810 2870
rect 6174 3346 6202 3351
rect 3840 2758 3972 2763
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3840 2725 3972 2730
rect 5996 2758 6128 2763
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 5996 2725 6128 2730
rect 2982 2647 2983 2673
rect 3009 2647 3010 2673
rect 2982 2641 3010 2647
rect 6174 2674 6202 3318
rect 6398 3345 6426 3351
rect 6398 3319 6399 3345
rect 6425 3319 6426 3345
rect 6398 3290 6426 3319
rect 6398 2842 6426 3262
rect 6510 3009 6538 3374
rect 6790 3369 6818 3374
rect 6734 3290 6762 3295
rect 6734 3243 6762 3262
rect 6846 3289 6874 4606
rect 6902 4241 6930 4774
rect 7074 4718 7206 4723
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7074 4685 7206 4690
rect 7238 4634 7266 4942
rect 6902 4215 6903 4241
rect 6929 4215 6930 4241
rect 6902 4209 6930 4215
rect 7070 4606 7266 4634
rect 7070 4073 7098 4606
rect 7294 4214 7322 5558
rect 7350 5194 7378 5199
rect 7350 4913 7378 5166
rect 7350 4887 7351 4913
rect 7377 4887 7378 4913
rect 7350 4881 7378 4887
rect 7070 4047 7071 4073
rect 7097 4047 7098 4073
rect 7070 4041 7098 4047
rect 7238 4186 7322 4214
rect 7406 4801 7434 4807
rect 7406 4775 7407 4801
rect 7433 4775 7434 4801
rect 7406 4186 7434 4775
rect 7462 4634 7490 4639
rect 7518 4634 7546 7238
rect 7574 7209 7602 7574
rect 8078 7569 8106 7574
rect 8152 7462 8284 7467
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8152 7429 8284 7434
rect 7574 7183 7575 7209
rect 7601 7183 7602 7209
rect 7574 7177 7602 7183
rect 7630 7209 7658 7215
rect 7630 7183 7631 7209
rect 7657 7183 7658 7209
rect 7630 6930 7658 7183
rect 8470 6986 8498 7911
rect 9230 7854 9362 7859
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9230 7821 9362 7826
rect 9230 7070 9362 7075
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9230 7037 9362 7042
rect 8470 6953 8498 6958
rect 7658 6902 7826 6930
rect 7630 6897 7658 6902
rect 7686 6706 7714 6711
rect 7574 6538 7602 6543
rect 7574 6482 7602 6510
rect 7574 6481 7658 6482
rect 7574 6455 7575 6481
rect 7601 6455 7658 6481
rect 7574 6454 7658 6455
rect 7574 6449 7602 6454
rect 7574 5978 7602 5983
rect 7574 5931 7602 5950
rect 7630 5810 7658 6454
rect 7686 6201 7714 6678
rect 7686 6175 7687 6201
rect 7713 6175 7714 6201
rect 7686 5922 7714 6175
rect 7742 5978 7770 5983
rect 7742 5931 7770 5950
rect 7686 5889 7714 5894
rect 7630 5782 7714 5810
rect 7490 4606 7546 4634
rect 7574 5754 7602 5759
rect 7602 5726 7658 5754
rect 7574 4913 7602 5726
rect 7630 5697 7658 5726
rect 7630 5671 7631 5697
rect 7657 5671 7658 5697
rect 7630 5665 7658 5671
rect 7686 5026 7714 5782
rect 7798 5698 7826 6902
rect 8152 6678 8284 6683
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8152 6645 8284 6650
rect 8974 6537 9002 6543
rect 8974 6511 8975 6537
rect 9001 6511 9002 6537
rect 7966 6482 7994 6487
rect 7966 6201 7994 6454
rect 7966 6175 7967 6201
rect 7993 6175 7994 6201
rect 7966 6169 7994 6175
rect 8022 6481 8050 6487
rect 8022 6455 8023 6481
rect 8049 6455 8050 6481
rect 8022 6145 8050 6455
rect 8974 6202 9002 6511
rect 9230 6286 9362 6291
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9230 6253 9362 6258
rect 8974 6169 9002 6174
rect 8022 6119 8023 6145
rect 8049 6119 8050 6145
rect 7686 4993 7714 4998
rect 7742 5670 7826 5698
rect 7910 6090 7938 6095
rect 7910 5977 7938 6062
rect 7910 5951 7911 5977
rect 7937 5951 7938 5977
rect 7742 4970 7770 5670
rect 7910 5642 7938 5951
rect 7742 4937 7770 4942
rect 7798 5614 7938 5642
rect 7966 5978 7994 5983
rect 7574 4887 7575 4913
rect 7601 4887 7602 4913
rect 7462 4601 7490 4606
rect 7574 4578 7602 4887
rect 7238 4018 7266 4186
rect 7406 4153 7434 4158
rect 7518 4577 7602 4578
rect 7518 4551 7575 4577
rect 7601 4551 7602 4577
rect 7518 4550 7602 4551
rect 7074 3934 7206 3939
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7074 3901 7206 3906
rect 7070 3850 7098 3855
rect 6958 3738 6986 3743
rect 6958 3691 6986 3710
rect 6846 3263 6847 3289
rect 6873 3263 6874 3289
rect 6510 2983 6511 3009
rect 6537 2983 6538 3009
rect 6510 2977 6538 2983
rect 6846 3234 6874 3263
rect 6398 2809 6426 2814
rect 6174 2641 6202 2646
rect 6846 2617 6874 3206
rect 7014 3626 7042 3631
rect 7014 3066 7042 3598
rect 7070 3289 7098 3822
rect 7182 3458 7210 3463
rect 7238 3458 7266 3990
rect 7518 4129 7546 4550
rect 7574 4545 7602 4550
rect 7798 4214 7826 5614
rect 7966 5586 7994 5950
rect 8022 5754 8050 6119
rect 8152 5894 8284 5899
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8152 5861 8284 5866
rect 8078 5754 8106 5759
rect 8022 5726 8078 5754
rect 8078 5721 8106 5726
rect 9086 5754 9114 5759
rect 9086 5707 9114 5726
rect 8022 5642 8050 5647
rect 8022 5595 8050 5614
rect 7910 5558 7994 5586
rect 7910 5305 7938 5558
rect 9230 5502 9362 5507
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9230 5469 9362 5474
rect 8134 5418 8162 5423
rect 7910 5279 7911 5305
rect 7937 5279 7938 5305
rect 7910 5273 7938 5279
rect 7966 5417 8162 5418
rect 7966 5391 8135 5417
rect 8161 5391 8162 5417
rect 7966 5390 8162 5391
rect 7910 4970 7938 4975
rect 7966 4970 7994 5390
rect 8134 5385 8162 5390
rect 8078 5306 8106 5311
rect 8078 5259 8106 5278
rect 8414 5306 8442 5311
rect 8694 5306 8722 5311
rect 8414 5305 8722 5306
rect 8414 5279 8415 5305
rect 8441 5279 8695 5305
rect 8721 5279 8722 5305
rect 8414 5278 8722 5279
rect 8414 5273 8442 5278
rect 8694 5273 8722 5278
rect 8302 5250 8330 5255
rect 8302 5249 8386 5250
rect 8302 5223 8303 5249
rect 8329 5223 8386 5249
rect 8302 5222 8386 5223
rect 8302 5217 8330 5222
rect 8190 5194 8218 5199
rect 8078 5193 8218 5194
rect 8078 5167 8191 5193
rect 8217 5167 8218 5193
rect 8078 5166 8218 5167
rect 8022 5026 8050 5031
rect 8078 5026 8106 5166
rect 8190 5161 8218 5166
rect 8152 5110 8284 5115
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8152 5077 8284 5082
rect 8050 4998 8106 5026
rect 8022 4993 8050 4998
rect 7910 4969 7994 4970
rect 7910 4943 7911 4969
rect 7937 4943 7994 4969
rect 7910 4942 7994 4943
rect 8302 4970 8330 4975
rect 8358 4970 8386 5222
rect 8330 4942 8386 4970
rect 8750 5249 8778 5255
rect 8750 5223 8751 5249
rect 8777 5223 8778 5249
rect 8750 4970 8778 5223
rect 8974 5249 9002 5255
rect 8974 5223 8975 5249
rect 9001 5223 9002 5249
rect 8918 5194 8946 5199
rect 8918 5147 8946 5166
rect 7910 4937 7938 4942
rect 8302 4937 8330 4942
rect 8750 4937 8778 4942
rect 8750 4578 8778 4583
rect 8750 4577 8834 4578
rect 8750 4551 8751 4577
rect 8777 4551 8834 4577
rect 8750 4550 8834 4551
rect 8750 4545 8778 4550
rect 8694 4521 8722 4527
rect 8694 4495 8695 4521
rect 8721 4495 8722 4521
rect 8152 4326 8284 4331
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8152 4293 8284 4298
rect 7518 4103 7519 4129
rect 7545 4103 7546 4129
rect 7210 3430 7266 3458
rect 7350 3737 7378 3743
rect 7350 3711 7351 3737
rect 7377 3711 7378 3737
rect 7182 3345 7210 3430
rect 7182 3319 7183 3345
rect 7209 3319 7210 3345
rect 7182 3313 7210 3319
rect 7070 3263 7071 3289
rect 7097 3263 7098 3289
rect 7070 3257 7098 3263
rect 7074 3150 7206 3155
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7074 3117 7206 3122
rect 7182 3066 7210 3071
rect 7014 3065 7210 3066
rect 7014 3039 7183 3065
rect 7209 3039 7210 3065
rect 7014 3038 7210 3039
rect 7182 3033 7210 3038
rect 7350 3010 7378 3711
rect 7518 3345 7546 4103
rect 7518 3319 7519 3345
rect 7545 3319 7546 3345
rect 7462 3066 7490 3071
rect 7462 3019 7490 3038
rect 6902 2954 6930 2959
rect 6902 2907 6930 2926
rect 7070 2898 7098 2903
rect 7070 2851 7098 2870
rect 7182 2898 7210 2903
rect 7182 2851 7210 2870
rect 7294 2674 7322 2679
rect 7294 2627 7322 2646
rect 6846 2591 6847 2617
rect 6873 2591 6874 2617
rect 6846 2585 6874 2591
rect 2926 2562 2954 2567
rect 2926 2515 2954 2534
rect 7350 2561 7378 2982
rect 7518 2954 7546 3319
rect 7742 4186 7826 4214
rect 7854 4186 7882 4191
rect 7742 3065 7770 4186
rect 7854 4139 7882 4158
rect 8302 3738 8330 3743
rect 7910 3682 7938 3687
rect 7910 3345 7938 3654
rect 8302 3681 8330 3710
rect 8302 3655 8303 3681
rect 8329 3655 8330 3681
rect 8302 3649 8330 3655
rect 8638 3737 8666 3743
rect 8638 3711 8639 3737
rect 8665 3711 8666 3737
rect 8152 3542 8284 3547
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8152 3509 8284 3514
rect 7910 3319 7911 3345
rect 7937 3319 7938 3345
rect 7910 3313 7938 3319
rect 8190 3346 8218 3351
rect 7742 3039 7743 3065
rect 7769 3039 7770 3065
rect 7742 3033 7770 3039
rect 8190 3066 8218 3318
rect 8134 3010 8162 3015
rect 8134 2963 8162 2982
rect 7518 2921 7546 2926
rect 7742 2954 7770 2959
rect 7742 2907 7770 2926
rect 8190 2953 8218 3038
rect 8190 2927 8191 2953
rect 8217 2927 8218 2953
rect 8190 2921 8218 2927
rect 8638 2954 8666 3711
rect 8694 3346 8722 4495
rect 8750 3682 8778 3687
rect 8750 3635 8778 3654
rect 8694 3313 8722 3318
rect 8806 3458 8834 4550
rect 8862 4521 8890 4527
rect 8862 4495 8863 4521
rect 8889 4495 8890 4521
rect 8862 3793 8890 4495
rect 8974 4214 9002 5223
rect 9030 4970 9058 4975
rect 9030 4923 9058 4942
rect 9230 4718 9362 4723
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9230 4685 9362 4690
rect 8862 3767 8863 3793
rect 8889 3767 8890 3793
rect 8862 3761 8890 3767
rect 8918 4186 9002 4214
rect 8918 4185 8946 4186
rect 8918 4159 8919 4185
rect 8945 4159 8946 4185
rect 8918 3794 8946 4159
rect 9230 3934 9362 3939
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9230 3901 9362 3906
rect 8918 3761 8946 3766
rect 8974 3738 9002 3743
rect 8974 3737 9058 3738
rect 8974 3711 8975 3737
rect 9001 3711 9058 3737
rect 8974 3710 9058 3711
rect 8974 3705 9002 3710
rect 8806 3430 9002 3458
rect 8750 3234 8778 3239
rect 8750 3065 8778 3206
rect 8750 3039 8751 3065
rect 8777 3039 8778 3065
rect 8750 3033 8778 3039
rect 8806 3010 8834 3430
rect 8974 3401 9002 3430
rect 8974 3375 8975 3401
rect 9001 3375 9002 3401
rect 8974 3369 9002 3375
rect 9030 3234 9058 3710
rect 9030 3201 9058 3206
rect 9230 3150 9362 3155
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9230 3117 9362 3122
rect 8806 2977 8834 2982
rect 8638 2921 8666 2926
rect 7406 2897 7434 2903
rect 7406 2871 7407 2897
rect 7433 2871 7434 2897
rect 7406 2842 7434 2871
rect 7406 2809 7434 2814
rect 8918 2842 8946 2847
rect 8152 2758 8284 2763
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8152 2725 8284 2730
rect 7350 2535 7351 2561
rect 7377 2535 7378 2561
rect 7350 2529 7378 2535
rect 2762 2366 2894 2371
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2762 2333 2894 2338
rect 4918 2366 5050 2371
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 4918 2333 5050 2338
rect 7074 2366 7206 2371
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7074 2333 7206 2338
rect 3840 1974 3972 1979
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3840 1941 3972 1946
rect 5996 1974 6128 1979
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 5996 1941 6128 1946
rect 8152 1974 8284 1979
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8152 1941 8284 1946
rect 2142 1777 2450 1778
rect 2142 1751 2143 1777
rect 2169 1751 2450 1777
rect 2142 1750 2450 1751
rect 2142 1745 2170 1750
rect 8806 1721 8834 1727
rect 8806 1695 8807 1721
rect 8833 1695 8834 1721
rect 8806 1666 8834 1695
rect 8918 1721 8946 2814
rect 9230 2366 9362 2371
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9230 2333 9362 2338
rect 8918 1695 8919 1721
rect 8945 1695 8946 1721
rect 8918 1689 8946 1695
rect 9086 1721 9114 1727
rect 9086 1695 9087 1721
rect 9113 1695 9114 1721
rect 8806 1633 8834 1638
rect 9086 1666 9114 1695
rect 2762 1582 2894 1587
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2762 1549 2894 1554
rect 4918 1582 5050 1587
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 4918 1549 5050 1554
rect 7074 1582 7206 1587
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7074 1549 7206 1554
rect 9086 1274 9114 1638
rect 9230 1582 9362 1587
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9230 1549 9362 1554
rect 9086 1241 9114 1246
rect 966 625 994 630
<< via2 >>
rect 1190 9198 1218 9226
rect 1684 8245 1712 8246
rect 1684 8219 1685 8245
rect 1685 8219 1711 8245
rect 1711 8219 1712 8245
rect 1684 8218 1712 8219
rect 1736 8245 1764 8246
rect 1736 8219 1737 8245
rect 1737 8219 1763 8245
rect 1763 8219 1764 8245
rect 1736 8218 1764 8219
rect 1788 8245 1816 8246
rect 1788 8219 1789 8245
rect 1789 8219 1815 8245
rect 1815 8219 1816 8245
rect 1788 8218 1816 8219
rect 854 7993 882 7994
rect 854 7967 855 7993
rect 855 7967 881 7993
rect 881 7967 882 7993
rect 854 7966 882 7967
rect 1078 7769 1106 7770
rect 1078 7743 1079 7769
rect 1079 7743 1105 7769
rect 1105 7743 1106 7769
rect 1078 7742 1106 7743
rect 1582 7993 1610 7994
rect 1582 7967 1583 7993
rect 1583 7967 1609 7993
rect 1609 7967 1610 7993
rect 1582 7966 1610 7967
rect 1190 7742 1218 7770
rect 1470 7657 1498 7658
rect 1470 7631 1471 7657
rect 1471 7631 1497 7657
rect 1497 7631 1498 7657
rect 1470 7630 1498 7631
rect 3840 8245 3868 8246
rect 3840 8219 3841 8245
rect 3841 8219 3867 8245
rect 3867 8219 3868 8245
rect 3840 8218 3868 8219
rect 3892 8245 3920 8246
rect 3892 8219 3893 8245
rect 3893 8219 3919 8245
rect 3919 8219 3920 8245
rect 3892 8218 3920 8219
rect 3944 8245 3972 8246
rect 3944 8219 3945 8245
rect 3945 8219 3971 8245
rect 3971 8219 3972 8245
rect 3944 8218 3972 8219
rect 5996 8245 6024 8246
rect 5996 8219 5997 8245
rect 5997 8219 6023 8245
rect 6023 8219 6024 8245
rect 5996 8218 6024 8219
rect 6048 8245 6076 8246
rect 6048 8219 6049 8245
rect 6049 8219 6075 8245
rect 6075 8219 6076 8245
rect 6048 8218 6076 8219
rect 6100 8245 6128 8246
rect 6100 8219 6101 8245
rect 6101 8219 6127 8245
rect 6127 8219 6128 8245
rect 6100 8218 6128 8219
rect 7462 8638 7490 8666
rect 8152 8245 8180 8246
rect 8152 8219 8153 8245
rect 8153 8219 8179 8245
rect 8179 8219 8180 8245
rect 8152 8218 8180 8219
rect 8204 8245 8232 8246
rect 8204 8219 8205 8245
rect 8205 8219 8231 8245
rect 8231 8219 8232 8245
rect 8204 8218 8232 8219
rect 8256 8245 8284 8246
rect 8256 8219 8257 8245
rect 8257 8219 8283 8245
rect 8283 8219 8284 8245
rect 8256 8218 8284 8219
rect 7406 8022 7434 8050
rect 2762 7853 2790 7854
rect 2762 7827 2763 7853
rect 2763 7827 2789 7853
rect 2789 7827 2790 7853
rect 2762 7826 2790 7827
rect 2814 7853 2842 7854
rect 2814 7827 2815 7853
rect 2815 7827 2841 7853
rect 2841 7827 2842 7853
rect 2814 7826 2842 7827
rect 2866 7853 2894 7854
rect 2866 7827 2867 7853
rect 2867 7827 2893 7853
rect 2893 7827 2894 7853
rect 2866 7826 2894 7827
rect 4918 7853 4946 7854
rect 4918 7827 4919 7853
rect 4919 7827 4945 7853
rect 4945 7827 4946 7853
rect 4918 7826 4946 7827
rect 4970 7853 4998 7854
rect 4970 7827 4971 7853
rect 4971 7827 4997 7853
rect 4997 7827 4998 7853
rect 4970 7826 4998 7827
rect 5022 7853 5050 7854
rect 5022 7827 5023 7853
rect 5023 7827 5049 7853
rect 5049 7827 5050 7853
rect 5022 7826 5050 7827
rect 7074 7853 7102 7854
rect 7074 7827 7075 7853
rect 7075 7827 7101 7853
rect 7101 7827 7102 7853
rect 7074 7826 7102 7827
rect 7126 7853 7154 7854
rect 7126 7827 7127 7853
rect 7127 7827 7153 7853
rect 7153 7827 7154 7853
rect 7126 7826 7154 7827
rect 7178 7853 7206 7854
rect 7178 7827 7179 7853
rect 7179 7827 7205 7853
rect 7205 7827 7206 7853
rect 7178 7826 7206 7827
rect 2870 7574 2898 7602
rect 3150 7630 3178 7658
rect 2478 7518 2506 7546
rect 1684 7461 1712 7462
rect 1684 7435 1685 7461
rect 1685 7435 1711 7461
rect 1711 7435 1712 7461
rect 1684 7434 1712 7435
rect 1736 7461 1764 7462
rect 1736 7435 1737 7461
rect 1737 7435 1763 7461
rect 1763 7435 1764 7461
rect 1736 7434 1764 7435
rect 1788 7461 1816 7462
rect 1788 7435 1789 7461
rect 1789 7435 1815 7461
rect 1815 7435 1816 7461
rect 1788 7434 1816 7435
rect 2982 7294 3010 7322
rect 854 6734 882 6762
rect 1246 6734 1274 6762
rect 1078 6174 1106 6202
rect 2762 7069 2790 7070
rect 2762 7043 2763 7069
rect 2763 7043 2789 7069
rect 2789 7043 2790 7069
rect 2762 7042 2790 7043
rect 2814 7069 2842 7070
rect 2814 7043 2815 7069
rect 2815 7043 2841 7069
rect 2841 7043 2842 7069
rect 2814 7042 2842 7043
rect 2866 7069 2894 7070
rect 2866 7043 2867 7069
rect 2867 7043 2893 7069
rect 2893 7043 2894 7069
rect 2866 7042 2894 7043
rect 2646 6958 2674 6986
rect 1684 6677 1712 6678
rect 1684 6651 1685 6677
rect 1685 6651 1711 6677
rect 1711 6651 1712 6677
rect 1684 6650 1712 6651
rect 1736 6677 1764 6678
rect 1736 6651 1737 6677
rect 1737 6651 1763 6677
rect 1763 6651 1764 6677
rect 1736 6650 1764 6651
rect 1788 6677 1816 6678
rect 1788 6651 1789 6677
rect 1789 6651 1815 6677
rect 1815 6651 1816 6677
rect 1788 6650 1816 6651
rect 4102 7574 4130 7602
rect 3840 7461 3868 7462
rect 3840 7435 3841 7461
rect 3841 7435 3867 7461
rect 3867 7435 3868 7461
rect 3840 7434 3868 7435
rect 3892 7461 3920 7462
rect 3892 7435 3893 7461
rect 3893 7435 3919 7461
rect 3919 7435 3920 7461
rect 3892 7434 3920 7435
rect 3944 7461 3972 7462
rect 3944 7435 3945 7461
rect 3945 7435 3971 7461
rect 3971 7435 3972 7461
rect 3944 7434 3972 7435
rect 3598 7321 3626 7322
rect 3598 7295 3599 7321
rect 3599 7295 3625 7321
rect 3625 7295 3626 7321
rect 3598 7294 3626 7295
rect 3766 7294 3794 7322
rect 3262 7265 3290 7266
rect 3262 7239 3263 7265
rect 3263 7239 3289 7265
rect 3289 7239 3290 7265
rect 3262 7238 3290 7239
rect 3318 7182 3346 7210
rect 1974 6174 2002 6202
rect 1582 6089 1610 6090
rect 1582 6063 1583 6089
rect 1583 6063 1609 6089
rect 1609 6063 1610 6089
rect 1582 6062 1610 6063
rect 2478 6174 2506 6202
rect 854 5502 882 5530
rect 1684 5893 1712 5894
rect 1684 5867 1685 5893
rect 1685 5867 1711 5893
rect 1711 5867 1712 5893
rect 1684 5866 1712 5867
rect 1736 5893 1764 5894
rect 1736 5867 1737 5893
rect 1737 5867 1763 5893
rect 1763 5867 1764 5893
rect 1736 5866 1764 5867
rect 1788 5893 1816 5894
rect 1788 5867 1789 5893
rect 1789 5867 1815 5893
rect 1815 5867 1816 5893
rect 1788 5866 1816 5867
rect 1190 5558 1218 5586
rect 2142 5558 2170 5586
rect 1134 5390 1162 5418
rect 1022 5222 1050 5250
rect 1246 5502 1274 5530
rect 1414 5249 1442 5250
rect 1414 5223 1415 5249
rect 1415 5223 1441 5249
rect 1441 5223 1442 5249
rect 1414 5222 1442 5223
rect 2366 5894 2394 5922
rect 2310 5361 2338 5362
rect 2310 5335 2311 5361
rect 2311 5335 2337 5361
rect 2337 5335 2338 5361
rect 2310 5334 2338 5335
rect 2198 5166 2226 5194
rect 1684 5109 1712 5110
rect 1684 5083 1685 5109
rect 1685 5083 1711 5109
rect 1711 5083 1712 5109
rect 1684 5082 1712 5083
rect 1736 5109 1764 5110
rect 1736 5083 1737 5109
rect 1737 5083 1763 5109
rect 1763 5083 1764 5109
rect 1736 5082 1764 5083
rect 1788 5109 1816 5110
rect 1788 5083 1789 5109
rect 1789 5083 1815 5109
rect 1815 5083 1816 5109
rect 1788 5082 1816 5083
rect 1470 4942 1498 4970
rect 1638 4998 1666 5026
rect 854 4270 882 4298
rect 1414 4550 1442 4578
rect 1526 4494 1554 4522
rect 1246 4270 1274 4298
rect 1470 4382 1498 4410
rect 2534 5894 2562 5922
rect 2478 5054 2506 5082
rect 1694 4942 1722 4970
rect 2590 5166 2618 5194
rect 2646 5361 2674 5362
rect 2646 5335 2647 5361
rect 2647 5335 2673 5361
rect 2673 5335 2674 5361
rect 2646 5334 2674 5335
rect 2646 5054 2674 5082
rect 2030 4830 2058 4858
rect 2534 4886 2562 4914
rect 2366 4550 2394 4578
rect 2142 4521 2170 4522
rect 2142 4495 2143 4521
rect 2143 4495 2169 4521
rect 2169 4495 2170 4521
rect 2142 4494 2170 4495
rect 2422 4830 2450 4858
rect 2086 4382 2114 4410
rect 2310 4409 2338 4410
rect 2310 4383 2311 4409
rect 2311 4383 2337 4409
rect 2337 4383 2338 4409
rect 2310 4382 2338 4383
rect 1684 4325 1712 4326
rect 1684 4299 1685 4325
rect 1685 4299 1711 4325
rect 1711 4299 1712 4325
rect 1684 4298 1712 4299
rect 1736 4325 1764 4326
rect 1736 4299 1737 4325
rect 1737 4299 1763 4325
rect 1763 4299 1764 4325
rect 1736 4298 1764 4299
rect 1788 4325 1816 4326
rect 1788 4299 1789 4325
rect 1789 4299 1815 4325
rect 1815 4299 1816 4325
rect 1788 4298 1816 4299
rect 2762 6285 2790 6286
rect 2762 6259 2763 6285
rect 2763 6259 2789 6285
rect 2789 6259 2790 6285
rect 2762 6258 2790 6259
rect 2814 6285 2842 6286
rect 2814 6259 2815 6285
rect 2815 6259 2841 6285
rect 2841 6259 2842 6285
rect 2814 6258 2842 6259
rect 2866 6285 2894 6286
rect 2866 6259 2867 6285
rect 2867 6259 2893 6285
rect 2893 6259 2894 6285
rect 2866 6258 2894 6259
rect 3654 7265 3682 7266
rect 3654 7239 3655 7265
rect 3655 7239 3681 7265
rect 3681 7239 3682 7265
rect 3654 7238 3682 7239
rect 4270 7294 4298 7322
rect 4438 7518 4466 7546
rect 3206 6958 3234 6986
rect 2982 6062 3010 6090
rect 2762 5501 2790 5502
rect 2762 5475 2763 5501
rect 2763 5475 2789 5501
rect 2789 5475 2790 5501
rect 2762 5474 2790 5475
rect 2814 5501 2842 5502
rect 2814 5475 2815 5501
rect 2815 5475 2841 5501
rect 2841 5475 2842 5501
rect 2814 5474 2842 5475
rect 2866 5501 2894 5502
rect 2866 5475 2867 5501
rect 2867 5475 2893 5501
rect 2893 5475 2894 5501
rect 2866 5474 2894 5475
rect 2814 5390 2842 5418
rect 2926 4857 2954 4858
rect 2926 4831 2927 4857
rect 2927 4831 2953 4857
rect 2953 4831 2954 4857
rect 2926 4830 2954 4831
rect 2762 4717 2790 4718
rect 2762 4691 2763 4717
rect 2763 4691 2789 4717
rect 2789 4691 2790 4717
rect 2762 4690 2790 4691
rect 2814 4717 2842 4718
rect 2814 4691 2815 4717
rect 2815 4691 2841 4717
rect 2841 4691 2842 4717
rect 2814 4690 2842 4691
rect 2866 4717 2894 4718
rect 2866 4691 2867 4717
rect 2867 4691 2893 4717
rect 2893 4691 2894 4717
rect 2866 4690 2894 4691
rect 3206 5110 3234 5138
rect 3150 5054 3178 5082
rect 2534 4494 2562 4522
rect 3542 6958 3570 6986
rect 3878 6958 3906 6986
rect 3990 6790 4018 6818
rect 3840 6677 3868 6678
rect 3840 6651 3841 6677
rect 3841 6651 3867 6677
rect 3867 6651 3868 6677
rect 3840 6650 3868 6651
rect 3892 6677 3920 6678
rect 3892 6651 3893 6677
rect 3893 6651 3919 6677
rect 3919 6651 3920 6677
rect 3892 6650 3920 6651
rect 3944 6677 3972 6678
rect 3944 6651 3945 6677
rect 3945 6651 3971 6677
rect 3971 6651 3972 6677
rect 3944 6650 3972 6651
rect 3654 6454 3682 6482
rect 3486 6174 3514 6202
rect 3318 6089 3346 6090
rect 3318 6063 3319 6089
rect 3319 6063 3345 6089
rect 3345 6063 3346 6089
rect 3318 6062 3346 6063
rect 3262 4942 3290 4970
rect 3318 5894 3346 5922
rect 3840 5893 3868 5894
rect 3840 5867 3841 5893
rect 3841 5867 3867 5893
rect 3867 5867 3868 5893
rect 3840 5866 3868 5867
rect 3892 5893 3920 5894
rect 3892 5867 3893 5893
rect 3893 5867 3919 5893
rect 3919 5867 3920 5893
rect 3892 5866 3920 5867
rect 3944 5893 3972 5894
rect 3944 5867 3945 5893
rect 3945 5867 3971 5893
rect 3971 5867 3972 5893
rect 3944 5866 3972 5867
rect 3374 5110 3402 5138
rect 3430 5390 3458 5418
rect 3318 4606 3346 4634
rect 3318 4521 3346 4522
rect 3318 4495 3319 4521
rect 3319 4495 3345 4521
rect 3345 4495 3346 4521
rect 3318 4494 3346 4495
rect 3206 4382 3234 4410
rect 2926 3990 2954 4018
rect 2762 3933 2790 3934
rect 2762 3907 2763 3933
rect 2763 3907 2789 3933
rect 2789 3907 2790 3933
rect 2762 3906 2790 3907
rect 2814 3933 2842 3934
rect 2814 3907 2815 3933
rect 2815 3907 2841 3933
rect 2841 3907 2842 3933
rect 2814 3906 2842 3907
rect 2866 3933 2894 3934
rect 2866 3907 2867 3933
rect 2867 3907 2893 3933
rect 2893 3907 2894 3933
rect 2866 3906 2894 3907
rect 2702 3849 2730 3850
rect 2702 3823 2703 3849
rect 2703 3823 2729 3849
rect 2729 3823 2730 3849
rect 2702 3822 2730 3823
rect 2982 3737 3010 3738
rect 2982 3711 2983 3737
rect 2983 3711 3009 3737
rect 3009 3711 3010 3737
rect 2982 3710 3010 3711
rect 1684 3541 1712 3542
rect 1684 3515 1685 3541
rect 1685 3515 1711 3541
rect 1711 3515 1712 3541
rect 1684 3514 1712 3515
rect 1736 3541 1764 3542
rect 1736 3515 1737 3541
rect 1737 3515 1763 3541
rect 1763 3515 1764 3541
rect 1736 3514 1764 3515
rect 1788 3541 1816 3542
rect 1788 3515 1789 3541
rect 1789 3515 1815 3541
rect 1815 3515 1816 3541
rect 1788 3514 1816 3515
rect 1470 3345 1498 3346
rect 1470 3319 1471 3345
rect 1471 3319 1497 3345
rect 1497 3319 1498 3345
rect 1470 3318 1498 3319
rect 854 3038 882 3066
rect 1246 3038 1274 3066
rect 1684 2757 1712 2758
rect 1684 2731 1685 2757
rect 1685 2731 1711 2757
rect 1711 2731 1712 2757
rect 1684 2730 1712 2731
rect 1736 2757 1764 2758
rect 1736 2731 1737 2757
rect 1737 2731 1763 2757
rect 1763 2731 1764 2757
rect 1736 2730 1764 2731
rect 1788 2757 1816 2758
rect 1788 2731 1789 2757
rect 1789 2731 1815 2757
rect 1815 2731 1816 2757
rect 1788 2730 1816 2731
rect 1022 2534 1050 2562
rect 854 2086 882 2114
rect 1246 2113 1274 2114
rect 1246 2087 1247 2113
rect 1247 2087 1273 2113
rect 1273 2087 1274 2113
rect 1246 2086 1274 2087
rect 1684 1973 1712 1974
rect 1684 1947 1685 1973
rect 1685 1947 1711 1973
rect 1711 1947 1712 1973
rect 1684 1946 1712 1947
rect 1736 1973 1764 1974
rect 1736 1947 1737 1973
rect 1737 1947 1763 1973
rect 1763 1947 1764 1973
rect 1736 1946 1764 1947
rect 1788 1973 1816 1974
rect 1788 1947 1789 1973
rect 1789 1947 1815 1973
rect 1815 1947 1816 1973
rect 1788 1946 1816 1947
rect 854 1806 882 1834
rect 2870 3598 2898 3626
rect 2762 3149 2790 3150
rect 2762 3123 2763 3149
rect 2763 3123 2789 3149
rect 2789 3123 2790 3149
rect 2762 3122 2790 3123
rect 2814 3149 2842 3150
rect 2814 3123 2815 3149
rect 2815 3123 2841 3149
rect 2841 3123 2842 3149
rect 2814 3122 2842 3123
rect 2866 3149 2894 3150
rect 2866 3123 2867 3149
rect 2867 3123 2893 3149
rect 2893 3123 2894 3149
rect 2866 3122 2894 3123
rect 4102 5390 4130 5418
rect 4158 6790 4186 6818
rect 3840 5109 3868 5110
rect 3840 5083 3841 5109
rect 3841 5083 3867 5109
rect 3867 5083 3868 5109
rect 3840 5082 3868 5083
rect 3892 5109 3920 5110
rect 3892 5083 3893 5109
rect 3893 5083 3919 5109
rect 3919 5083 3920 5109
rect 3892 5082 3920 5083
rect 3944 5109 3972 5110
rect 3944 5083 3945 5109
rect 3945 5083 3971 5109
rect 3971 5083 3972 5109
rect 3944 5082 3972 5083
rect 3542 4969 3570 4970
rect 3542 4943 3543 4969
rect 3543 4943 3569 4969
rect 3569 4943 3570 4969
rect 3542 4942 3570 4943
rect 4046 4801 4074 4802
rect 4046 4775 4047 4801
rect 4047 4775 4073 4801
rect 4073 4775 4074 4801
rect 4046 4774 4074 4775
rect 3840 4325 3868 4326
rect 3840 4299 3841 4325
rect 3841 4299 3867 4325
rect 3867 4299 3868 4325
rect 3840 4298 3868 4299
rect 3892 4325 3920 4326
rect 3892 4299 3893 4325
rect 3893 4299 3919 4325
rect 3919 4299 3920 4325
rect 3892 4298 3920 4299
rect 3944 4325 3972 4326
rect 3944 4299 3945 4325
rect 3945 4299 3971 4325
rect 3971 4299 3972 4325
rect 3944 4298 3972 4299
rect 3822 4214 3850 4242
rect 3374 3849 3402 3850
rect 3374 3823 3375 3849
rect 3375 3823 3401 3849
rect 3401 3823 3402 3849
rect 3374 3822 3402 3823
rect 3206 3766 3234 3794
rect 3318 3737 3346 3738
rect 3318 3711 3319 3737
rect 3319 3711 3345 3737
rect 3345 3711 3346 3737
rect 3318 3710 3346 3711
rect 4214 6174 4242 6202
rect 4382 6089 4410 6090
rect 4382 6063 4383 6089
rect 4383 6063 4409 6089
rect 4409 6063 4410 6089
rect 4382 6062 4410 6063
rect 4494 7209 4522 7210
rect 4494 7183 4495 7209
rect 4495 7183 4521 7209
rect 4521 7183 4522 7209
rect 4494 7182 4522 7183
rect 4942 7126 4970 7154
rect 5110 7182 5138 7210
rect 4918 7069 4946 7070
rect 4918 7043 4919 7069
rect 4919 7043 4945 7069
rect 4945 7043 4946 7069
rect 4918 7042 4946 7043
rect 4970 7069 4998 7070
rect 4970 7043 4971 7069
rect 4971 7043 4997 7069
rect 4997 7043 4998 7069
rect 4970 7042 4998 7043
rect 5022 7069 5050 7070
rect 5022 7043 5023 7069
rect 5023 7043 5049 7069
rect 5049 7043 5050 7069
rect 5022 7042 5050 7043
rect 4494 6201 4522 6202
rect 4494 6175 4495 6201
rect 4495 6175 4521 6201
rect 4521 6175 4522 6201
rect 4494 6174 4522 6175
rect 4662 6369 4690 6370
rect 4662 6343 4663 6369
rect 4663 6343 4689 6369
rect 4689 6343 4690 6369
rect 4662 6342 4690 6343
rect 5166 6846 5194 6874
rect 5054 6425 5082 6426
rect 5054 6399 5055 6425
rect 5055 6399 5081 6425
rect 5081 6399 5082 6425
rect 5054 6398 5082 6399
rect 4918 6285 4946 6286
rect 4918 6259 4919 6285
rect 4919 6259 4945 6285
rect 4945 6259 4946 6285
rect 4918 6258 4946 6259
rect 4970 6285 4998 6286
rect 4970 6259 4971 6285
rect 4971 6259 4997 6285
rect 4997 6259 4998 6285
rect 4970 6258 4998 6259
rect 5022 6285 5050 6286
rect 5022 6259 5023 6285
rect 5023 6259 5049 6285
rect 5049 6259 5050 6285
rect 5022 6258 5050 6259
rect 4830 6201 4858 6202
rect 4830 6175 4831 6201
rect 4831 6175 4857 6201
rect 4857 6175 4858 6201
rect 4830 6174 4858 6175
rect 4550 6118 4578 6146
rect 4886 6118 4914 6146
rect 4942 6089 4970 6090
rect 4942 6063 4943 6089
rect 4943 6063 4969 6089
rect 4969 6063 4970 6089
rect 4942 6062 4970 6063
rect 5110 6006 5138 6034
rect 4550 5558 4578 5586
rect 4494 5417 4522 5418
rect 4494 5391 4495 5417
rect 4495 5391 4521 5417
rect 4521 5391 4522 5417
rect 4494 5390 4522 5391
rect 5334 6790 5362 6818
rect 5614 6929 5642 6930
rect 5614 6903 5615 6929
rect 5615 6903 5641 6929
rect 5641 6903 5642 6929
rect 5614 6902 5642 6903
rect 5996 7461 6024 7462
rect 5996 7435 5997 7461
rect 5997 7435 6023 7461
rect 6023 7435 6024 7461
rect 5996 7434 6024 7435
rect 6048 7461 6076 7462
rect 6048 7435 6049 7461
rect 6049 7435 6075 7461
rect 6075 7435 6076 7461
rect 6048 7434 6076 7435
rect 6100 7461 6128 7462
rect 6100 7435 6101 7461
rect 6101 7435 6127 7461
rect 6127 7435 6128 7461
rect 6100 7434 6128 7435
rect 6174 7294 6202 7322
rect 5838 7070 5866 7098
rect 5894 6734 5922 6762
rect 6510 7070 6538 7098
rect 6118 6873 6146 6874
rect 6118 6847 6119 6873
rect 6119 6847 6145 6873
rect 6145 6847 6146 6873
rect 6118 6846 6146 6847
rect 5996 6677 6024 6678
rect 5996 6651 5997 6677
rect 5997 6651 6023 6677
rect 6023 6651 6024 6677
rect 5996 6650 6024 6651
rect 6048 6677 6076 6678
rect 6048 6651 6049 6677
rect 6049 6651 6075 6677
rect 6075 6651 6076 6677
rect 6048 6650 6076 6651
rect 6100 6677 6128 6678
rect 6100 6651 6101 6677
rect 6101 6651 6127 6677
rect 6127 6651 6128 6677
rect 6100 6650 6128 6651
rect 6174 6566 6202 6594
rect 5222 6145 5250 6146
rect 5222 6119 5223 6145
rect 5223 6119 5249 6145
rect 5249 6119 5250 6145
rect 5222 6118 5250 6119
rect 5334 5894 5362 5922
rect 4918 5501 4946 5502
rect 4918 5475 4919 5501
rect 4919 5475 4945 5501
rect 4945 5475 4946 5501
rect 4918 5474 4946 5475
rect 4970 5501 4998 5502
rect 4970 5475 4971 5501
rect 4971 5475 4997 5501
rect 4997 5475 4998 5501
rect 4970 5474 4998 5475
rect 5022 5501 5050 5502
rect 5022 5475 5023 5501
rect 5023 5475 5049 5501
rect 5049 5475 5050 5501
rect 5022 5474 5050 5475
rect 5222 5558 5250 5586
rect 4326 4942 4354 4970
rect 4830 5249 4858 5250
rect 4830 5223 4831 5249
rect 4831 5223 4857 5249
rect 4857 5223 4858 5249
rect 4830 5222 4858 5223
rect 4718 5166 4746 5194
rect 4382 4774 4410 4802
rect 4438 4718 4466 4746
rect 4494 4774 4522 4802
rect 4158 3990 4186 4018
rect 4214 4438 4242 4466
rect 3430 3598 3458 3626
rect 3878 3737 3906 3738
rect 3878 3711 3879 3737
rect 3879 3711 3905 3737
rect 3905 3711 3906 3737
rect 3878 3710 3906 3711
rect 4326 4521 4354 4522
rect 4326 4495 4327 4521
rect 4327 4495 4353 4521
rect 4353 4495 4354 4521
rect 4326 4494 4354 4495
rect 4550 4550 4578 4578
rect 4494 4494 4522 4522
rect 4830 4913 4858 4914
rect 4830 4887 4831 4913
rect 4831 4887 4857 4913
rect 4857 4887 4858 4913
rect 4830 4886 4858 4887
rect 4774 4857 4802 4858
rect 4774 4831 4775 4857
rect 4775 4831 4801 4857
rect 4801 4831 4802 4857
rect 4774 4830 4802 4831
rect 4830 4718 4858 4746
rect 4918 4717 4946 4718
rect 4918 4691 4919 4717
rect 4919 4691 4945 4717
rect 4945 4691 4946 4717
rect 4918 4690 4946 4691
rect 4970 4717 4998 4718
rect 4970 4691 4971 4717
rect 4971 4691 4997 4717
rect 4997 4691 4998 4717
rect 4970 4690 4998 4691
rect 5022 4717 5050 4718
rect 5022 4691 5023 4717
rect 5023 4691 5049 4717
rect 5049 4691 5050 4717
rect 5022 4690 5050 4691
rect 5166 5390 5194 5418
rect 4830 4521 4858 4522
rect 4830 4495 4831 4521
rect 4831 4495 4857 4521
rect 4857 4495 4858 4521
rect 4830 4494 4858 4495
rect 5054 4270 5082 4298
rect 4270 4158 4298 4186
rect 4886 4185 4914 4186
rect 4886 4159 4887 4185
rect 4887 4159 4913 4185
rect 4913 4159 4914 4185
rect 4886 4158 4914 4159
rect 5446 4913 5474 4914
rect 5446 4887 5447 4913
rect 5447 4887 5473 4913
rect 5473 4887 5474 4913
rect 5446 4886 5474 4887
rect 5278 4830 5306 4858
rect 5502 4606 5530 4634
rect 5110 4102 5138 4130
rect 4918 3933 4946 3934
rect 4918 3907 4919 3933
rect 4919 3907 4945 3933
rect 4945 3907 4946 3933
rect 4918 3906 4946 3907
rect 4970 3933 4998 3934
rect 4970 3907 4971 3933
rect 4971 3907 4997 3933
rect 4997 3907 4998 3933
rect 4970 3906 4998 3907
rect 5022 3933 5050 3934
rect 5022 3907 5023 3933
rect 5023 3907 5049 3933
rect 5049 3907 5050 3933
rect 5022 3906 5050 3907
rect 4494 3849 4522 3850
rect 4494 3823 4495 3849
rect 4495 3823 4521 3849
rect 4521 3823 4522 3849
rect 4494 3822 4522 3823
rect 3766 3598 3794 3626
rect 4270 3598 4298 3626
rect 3840 3541 3868 3542
rect 3840 3515 3841 3541
rect 3841 3515 3867 3541
rect 3867 3515 3868 3541
rect 3840 3514 3868 3515
rect 3892 3541 3920 3542
rect 3892 3515 3893 3541
rect 3893 3515 3919 3541
rect 3919 3515 3920 3541
rect 3892 3514 3920 3515
rect 3944 3541 3972 3542
rect 3944 3515 3945 3541
rect 3945 3515 3971 3541
rect 3971 3515 3972 3541
rect 3944 3514 3972 3515
rect 3038 3318 3066 3346
rect 5110 3849 5138 3850
rect 5110 3823 5111 3849
rect 5111 3823 5137 3849
rect 5137 3823 5138 3849
rect 5110 3822 5138 3823
rect 4718 3793 4746 3794
rect 4718 3767 4719 3793
rect 4719 3767 4745 3793
rect 4745 3767 4746 3793
rect 4718 3766 4746 3767
rect 5334 4214 5362 4242
rect 5614 6174 5642 6202
rect 5838 6174 5866 6202
rect 5950 6286 5978 6314
rect 5670 6006 5698 6034
rect 6342 6342 6370 6370
rect 6006 6145 6034 6146
rect 6006 6119 6007 6145
rect 6007 6119 6033 6145
rect 6033 6119 6034 6145
rect 6006 6118 6034 6119
rect 6062 6089 6090 6090
rect 6062 6063 6063 6089
rect 6063 6063 6089 6089
rect 6089 6063 6090 6089
rect 6062 6062 6090 6063
rect 6230 6089 6258 6090
rect 6230 6063 6231 6089
rect 6231 6063 6257 6089
rect 6257 6063 6258 6089
rect 6230 6062 6258 6063
rect 5894 5894 5922 5922
rect 5838 5334 5866 5362
rect 5996 5893 6024 5894
rect 5996 5867 5997 5893
rect 5997 5867 6023 5893
rect 6023 5867 6024 5893
rect 5996 5866 6024 5867
rect 6048 5893 6076 5894
rect 6048 5867 6049 5893
rect 6049 5867 6075 5893
rect 6075 5867 6076 5893
rect 6048 5866 6076 5867
rect 6100 5893 6128 5894
rect 6100 5867 6101 5893
rect 6101 5867 6127 5893
rect 6127 5867 6128 5893
rect 6100 5866 6128 5867
rect 6174 5361 6202 5362
rect 6174 5335 6175 5361
rect 6175 5335 6201 5361
rect 6201 5335 6202 5361
rect 6174 5334 6202 5335
rect 5996 5109 6024 5110
rect 5996 5083 5997 5109
rect 5997 5083 6023 5109
rect 6023 5083 6024 5109
rect 5996 5082 6024 5083
rect 6048 5109 6076 5110
rect 6048 5083 6049 5109
rect 6049 5083 6075 5109
rect 6075 5083 6076 5109
rect 6048 5082 6076 5083
rect 6100 5109 6128 5110
rect 6100 5083 6101 5109
rect 6101 5083 6127 5109
rect 6127 5083 6128 5109
rect 6100 5082 6128 5083
rect 5894 4550 5922 4578
rect 6174 4550 6202 4578
rect 6342 5222 6370 5250
rect 5726 4270 5754 4298
rect 5222 4158 5250 4186
rect 5670 4158 5698 4186
rect 5334 4046 5362 4074
rect 5558 4129 5586 4130
rect 5558 4103 5559 4129
rect 5559 4103 5585 4129
rect 5585 4103 5586 4129
rect 5558 4102 5586 4103
rect 5558 3766 5586 3794
rect 4886 3737 4914 3738
rect 4886 3711 4887 3737
rect 4887 3711 4913 3737
rect 4913 3711 4914 3737
rect 4886 3710 4914 3711
rect 4830 3598 4858 3626
rect 4998 3345 5026 3346
rect 4998 3319 4999 3345
rect 4999 3319 5025 3345
rect 5025 3319 5026 3345
rect 4998 3318 5026 3319
rect 5222 3262 5250 3290
rect 4918 3149 4946 3150
rect 4918 3123 4919 3149
rect 4919 3123 4945 3149
rect 4945 3123 4946 3149
rect 4918 3122 4946 3123
rect 4970 3149 4998 3150
rect 4970 3123 4971 3149
rect 4971 3123 4997 3149
rect 4997 3123 4998 3149
rect 4970 3122 4998 3123
rect 5022 3149 5050 3150
rect 5022 3123 5023 3149
rect 5023 3123 5049 3149
rect 5049 3123 5050 3149
rect 5022 3122 5050 3123
rect 5996 4325 6024 4326
rect 5996 4299 5997 4325
rect 5997 4299 6023 4325
rect 6023 4299 6024 4325
rect 5996 4298 6024 4299
rect 6048 4325 6076 4326
rect 6048 4299 6049 4325
rect 6049 4299 6075 4325
rect 6075 4299 6076 4325
rect 6048 4298 6076 4299
rect 6100 4325 6128 4326
rect 6100 4299 6101 4325
rect 6101 4299 6127 4325
rect 6127 4299 6128 4325
rect 6100 4298 6128 4299
rect 6398 5614 6426 5642
rect 6454 4998 6482 5026
rect 8358 8022 8386 8050
rect 8582 8049 8610 8050
rect 8582 8023 8583 8049
rect 8583 8023 8609 8049
rect 8609 8023 8610 8049
rect 8582 8022 8610 8023
rect 6958 7265 6986 7266
rect 6958 7239 6959 7265
rect 6959 7239 6985 7265
rect 6985 7239 6986 7265
rect 6958 7238 6986 7239
rect 7074 7069 7102 7070
rect 7074 7043 7075 7069
rect 7075 7043 7101 7069
rect 7101 7043 7102 7069
rect 7074 7042 7102 7043
rect 7126 7069 7154 7070
rect 7126 7043 7127 7069
rect 7127 7043 7153 7069
rect 7153 7043 7154 7069
rect 7126 7042 7154 7043
rect 7178 7069 7206 7070
rect 7178 7043 7179 7069
rect 7179 7043 7205 7069
rect 7205 7043 7206 7069
rect 7178 7042 7206 7043
rect 7518 7238 7546 7266
rect 6790 6593 6818 6594
rect 6790 6567 6791 6593
rect 6791 6567 6817 6593
rect 6817 6567 6818 6593
rect 6790 6566 6818 6567
rect 6566 5726 6594 5754
rect 6622 6342 6650 6370
rect 6846 6369 6874 6370
rect 6846 6343 6847 6369
rect 6847 6343 6873 6369
rect 6873 6343 6874 6369
rect 6846 6342 6874 6343
rect 6902 6286 6930 6314
rect 6734 6118 6762 6146
rect 6846 6089 6874 6090
rect 6846 6063 6847 6089
rect 6847 6063 6873 6089
rect 6873 6063 6874 6089
rect 6846 6062 6874 6063
rect 6678 5977 6706 5978
rect 6678 5951 6679 5977
rect 6679 5951 6705 5977
rect 6705 5951 6706 5977
rect 6678 5950 6706 5951
rect 7462 6481 7490 6482
rect 7462 6455 7463 6481
rect 7463 6455 7489 6481
rect 7489 6455 7490 6481
rect 7462 6454 7490 6455
rect 7238 6342 7266 6370
rect 7074 6285 7102 6286
rect 7074 6259 7075 6285
rect 7075 6259 7101 6285
rect 7101 6259 7102 6285
rect 7074 6258 7102 6259
rect 7126 6285 7154 6286
rect 7126 6259 7127 6285
rect 7127 6259 7153 6285
rect 7153 6259 7154 6285
rect 7126 6258 7154 6259
rect 7178 6285 7206 6286
rect 7178 6259 7179 6285
rect 7179 6259 7205 6285
rect 7205 6259 7206 6285
rect 7178 6258 7206 6259
rect 7014 6174 7042 6202
rect 7238 6201 7266 6202
rect 7238 6175 7239 6201
rect 7239 6175 7265 6201
rect 7265 6175 7266 6201
rect 7238 6174 7266 6175
rect 6958 6062 6986 6090
rect 7406 6089 7434 6090
rect 7406 6063 7407 6089
rect 7407 6063 7433 6089
rect 7433 6063 7434 6089
rect 7406 6062 7434 6063
rect 6622 5670 6650 5698
rect 6510 4942 6538 4970
rect 6790 5782 6818 5810
rect 6734 4942 6762 4970
rect 6846 5697 6874 5698
rect 6846 5671 6847 5697
rect 6847 5671 6873 5697
rect 6873 5671 6874 5697
rect 6846 5670 6874 5671
rect 7126 5641 7154 5642
rect 7126 5615 7127 5641
rect 7127 5615 7153 5641
rect 7153 5615 7154 5641
rect 7126 5614 7154 5615
rect 7462 5614 7490 5642
rect 6958 5502 6986 5530
rect 7182 5585 7210 5586
rect 7182 5559 7183 5585
rect 7183 5559 7209 5585
rect 7209 5559 7210 5585
rect 7182 5558 7210 5559
rect 7074 5501 7102 5502
rect 7074 5475 7075 5501
rect 7075 5475 7101 5501
rect 7101 5475 7102 5501
rect 7074 5474 7102 5475
rect 7126 5501 7154 5502
rect 7126 5475 7127 5501
rect 7127 5475 7153 5501
rect 7153 5475 7154 5501
rect 7126 5474 7154 5475
rect 7178 5501 7206 5502
rect 7178 5475 7179 5501
rect 7179 5475 7205 5501
rect 7205 5475 7206 5501
rect 7178 5474 7206 5475
rect 7014 5278 7042 5306
rect 7014 4998 7042 5026
rect 7126 5025 7154 5026
rect 7126 4999 7127 5025
rect 7127 4999 7153 5025
rect 7153 4999 7154 5025
rect 7126 4998 7154 4999
rect 7238 4969 7266 4970
rect 7238 4943 7239 4969
rect 7239 4943 7265 4969
rect 7265 4943 7266 4969
rect 7238 4942 7266 4943
rect 6678 4774 6706 4802
rect 5894 4158 5922 4186
rect 6230 4129 6258 4130
rect 6230 4103 6231 4129
rect 6231 4103 6257 4129
rect 6257 4103 6258 4129
rect 6230 4102 6258 4103
rect 6622 4158 6650 4186
rect 6454 4129 6482 4130
rect 6454 4103 6455 4129
rect 6455 4103 6481 4129
rect 6481 4103 6482 4129
rect 6454 4102 6482 4103
rect 5894 4073 5922 4074
rect 5894 4047 5895 4073
rect 5895 4047 5921 4073
rect 5921 4047 5922 4073
rect 5894 4046 5922 4047
rect 6174 3822 6202 3850
rect 5838 3598 5866 3626
rect 5996 3541 6024 3542
rect 5996 3515 5997 3541
rect 5997 3515 6023 3541
rect 6023 3515 6024 3541
rect 5996 3514 6024 3515
rect 6048 3541 6076 3542
rect 6048 3515 6049 3541
rect 6049 3515 6075 3541
rect 6075 3515 6076 3541
rect 6048 3514 6076 3515
rect 6100 3541 6128 3542
rect 6100 3515 6101 3541
rect 6101 3515 6127 3541
rect 6127 3515 6128 3541
rect 6100 3514 6128 3515
rect 6230 3457 6258 3458
rect 6230 3431 6231 3457
rect 6231 3431 6257 3457
rect 6257 3431 6258 3457
rect 6230 3430 6258 3431
rect 6902 4774 6930 4802
rect 6846 4606 6874 4634
rect 6790 4102 6818 4130
rect 6790 3934 6818 3962
rect 6734 3822 6762 3850
rect 6286 3374 6314 3402
rect 5782 2870 5810 2898
rect 6174 3345 6202 3346
rect 6174 3319 6175 3345
rect 6175 3319 6201 3345
rect 6201 3319 6202 3345
rect 6174 3318 6202 3319
rect 3840 2757 3868 2758
rect 3840 2731 3841 2757
rect 3841 2731 3867 2757
rect 3867 2731 3868 2757
rect 3840 2730 3868 2731
rect 3892 2757 3920 2758
rect 3892 2731 3893 2757
rect 3893 2731 3919 2757
rect 3919 2731 3920 2757
rect 3892 2730 3920 2731
rect 3944 2757 3972 2758
rect 3944 2731 3945 2757
rect 3945 2731 3971 2757
rect 3971 2731 3972 2757
rect 3944 2730 3972 2731
rect 5996 2757 6024 2758
rect 5996 2731 5997 2757
rect 5997 2731 6023 2757
rect 6023 2731 6024 2757
rect 5996 2730 6024 2731
rect 6048 2757 6076 2758
rect 6048 2731 6049 2757
rect 6049 2731 6075 2757
rect 6075 2731 6076 2757
rect 6048 2730 6076 2731
rect 6100 2757 6128 2758
rect 6100 2731 6101 2757
rect 6101 2731 6127 2757
rect 6127 2731 6128 2757
rect 6100 2730 6128 2731
rect 6398 3262 6426 3290
rect 6734 3289 6762 3290
rect 6734 3263 6735 3289
rect 6735 3263 6761 3289
rect 6761 3263 6762 3289
rect 6734 3262 6762 3263
rect 7074 4717 7102 4718
rect 7074 4691 7075 4717
rect 7075 4691 7101 4717
rect 7101 4691 7102 4717
rect 7074 4690 7102 4691
rect 7126 4717 7154 4718
rect 7126 4691 7127 4717
rect 7127 4691 7153 4717
rect 7153 4691 7154 4717
rect 7126 4690 7154 4691
rect 7178 4717 7206 4718
rect 7178 4691 7179 4717
rect 7179 4691 7205 4717
rect 7205 4691 7206 4717
rect 7178 4690 7206 4691
rect 7350 5166 7378 5194
rect 8152 7461 8180 7462
rect 8152 7435 8153 7461
rect 8153 7435 8179 7461
rect 8179 7435 8180 7461
rect 8152 7434 8180 7435
rect 8204 7461 8232 7462
rect 8204 7435 8205 7461
rect 8205 7435 8231 7461
rect 8231 7435 8232 7461
rect 8204 7434 8232 7435
rect 8256 7461 8284 7462
rect 8256 7435 8257 7461
rect 8257 7435 8283 7461
rect 8283 7435 8284 7461
rect 8256 7434 8284 7435
rect 9230 7853 9258 7854
rect 9230 7827 9231 7853
rect 9231 7827 9257 7853
rect 9257 7827 9258 7853
rect 9230 7826 9258 7827
rect 9282 7853 9310 7854
rect 9282 7827 9283 7853
rect 9283 7827 9309 7853
rect 9309 7827 9310 7853
rect 9282 7826 9310 7827
rect 9334 7853 9362 7854
rect 9334 7827 9335 7853
rect 9335 7827 9361 7853
rect 9361 7827 9362 7853
rect 9334 7826 9362 7827
rect 9230 7069 9258 7070
rect 9230 7043 9231 7069
rect 9231 7043 9257 7069
rect 9257 7043 9258 7069
rect 9230 7042 9258 7043
rect 9282 7069 9310 7070
rect 9282 7043 9283 7069
rect 9283 7043 9309 7069
rect 9309 7043 9310 7069
rect 9282 7042 9310 7043
rect 9334 7069 9362 7070
rect 9334 7043 9335 7069
rect 9335 7043 9361 7069
rect 9361 7043 9362 7069
rect 9334 7042 9362 7043
rect 8470 6958 8498 6986
rect 7630 6902 7658 6930
rect 7686 6678 7714 6706
rect 7574 6510 7602 6538
rect 7574 5977 7602 5978
rect 7574 5951 7575 5977
rect 7575 5951 7601 5977
rect 7601 5951 7602 5977
rect 7574 5950 7602 5951
rect 7742 5977 7770 5978
rect 7742 5951 7743 5977
rect 7743 5951 7769 5977
rect 7769 5951 7770 5977
rect 7742 5950 7770 5951
rect 7686 5894 7714 5922
rect 7462 4606 7490 4634
rect 7574 5726 7602 5754
rect 8152 6677 8180 6678
rect 8152 6651 8153 6677
rect 8153 6651 8179 6677
rect 8179 6651 8180 6677
rect 8152 6650 8180 6651
rect 8204 6677 8232 6678
rect 8204 6651 8205 6677
rect 8205 6651 8231 6677
rect 8231 6651 8232 6677
rect 8204 6650 8232 6651
rect 8256 6677 8284 6678
rect 8256 6651 8257 6677
rect 8257 6651 8283 6677
rect 8283 6651 8284 6677
rect 8256 6650 8284 6651
rect 7966 6454 7994 6482
rect 9230 6285 9258 6286
rect 9230 6259 9231 6285
rect 9231 6259 9257 6285
rect 9257 6259 9258 6285
rect 9230 6258 9258 6259
rect 9282 6285 9310 6286
rect 9282 6259 9283 6285
rect 9283 6259 9309 6285
rect 9309 6259 9310 6285
rect 9282 6258 9310 6259
rect 9334 6285 9362 6286
rect 9334 6259 9335 6285
rect 9335 6259 9361 6285
rect 9361 6259 9362 6285
rect 9334 6258 9362 6259
rect 8974 6174 9002 6202
rect 7686 4998 7714 5026
rect 7910 6062 7938 6090
rect 7742 4942 7770 4970
rect 7966 5950 7994 5978
rect 7406 4158 7434 4186
rect 7238 4017 7266 4018
rect 7238 3991 7239 4017
rect 7239 3991 7265 4017
rect 7265 3991 7266 4017
rect 7238 3990 7266 3991
rect 7074 3933 7102 3934
rect 7074 3907 7075 3933
rect 7075 3907 7101 3933
rect 7101 3907 7102 3933
rect 7074 3906 7102 3907
rect 7126 3933 7154 3934
rect 7126 3907 7127 3933
rect 7127 3907 7153 3933
rect 7153 3907 7154 3933
rect 7126 3906 7154 3907
rect 7178 3933 7206 3934
rect 7178 3907 7179 3933
rect 7179 3907 7205 3933
rect 7205 3907 7206 3933
rect 7178 3906 7206 3907
rect 7070 3822 7098 3850
rect 6958 3737 6986 3738
rect 6958 3711 6959 3737
rect 6959 3711 6985 3737
rect 6985 3711 6986 3737
rect 6958 3710 6986 3711
rect 6846 3206 6874 3234
rect 6398 2814 6426 2842
rect 6174 2646 6202 2674
rect 7014 3598 7042 3626
rect 8152 5893 8180 5894
rect 8152 5867 8153 5893
rect 8153 5867 8179 5893
rect 8179 5867 8180 5893
rect 8152 5866 8180 5867
rect 8204 5893 8232 5894
rect 8204 5867 8205 5893
rect 8205 5867 8231 5893
rect 8231 5867 8232 5893
rect 8204 5866 8232 5867
rect 8256 5893 8284 5894
rect 8256 5867 8257 5893
rect 8257 5867 8283 5893
rect 8283 5867 8284 5893
rect 8256 5866 8284 5867
rect 8078 5726 8106 5754
rect 9086 5753 9114 5754
rect 9086 5727 9087 5753
rect 9087 5727 9113 5753
rect 9113 5727 9114 5753
rect 9086 5726 9114 5727
rect 8022 5641 8050 5642
rect 8022 5615 8023 5641
rect 8023 5615 8049 5641
rect 8049 5615 8050 5641
rect 8022 5614 8050 5615
rect 9230 5501 9258 5502
rect 9230 5475 9231 5501
rect 9231 5475 9257 5501
rect 9257 5475 9258 5501
rect 9230 5474 9258 5475
rect 9282 5501 9310 5502
rect 9282 5475 9283 5501
rect 9283 5475 9309 5501
rect 9309 5475 9310 5501
rect 9282 5474 9310 5475
rect 9334 5501 9362 5502
rect 9334 5475 9335 5501
rect 9335 5475 9361 5501
rect 9361 5475 9362 5501
rect 9334 5474 9362 5475
rect 8078 5305 8106 5306
rect 8078 5279 8079 5305
rect 8079 5279 8105 5305
rect 8105 5279 8106 5305
rect 8078 5278 8106 5279
rect 8152 5109 8180 5110
rect 8152 5083 8153 5109
rect 8153 5083 8179 5109
rect 8179 5083 8180 5109
rect 8152 5082 8180 5083
rect 8204 5109 8232 5110
rect 8204 5083 8205 5109
rect 8205 5083 8231 5109
rect 8231 5083 8232 5109
rect 8204 5082 8232 5083
rect 8256 5109 8284 5110
rect 8256 5083 8257 5109
rect 8257 5083 8283 5109
rect 8283 5083 8284 5109
rect 8256 5082 8284 5083
rect 8022 4998 8050 5026
rect 8302 4942 8330 4970
rect 8918 5193 8946 5194
rect 8918 5167 8919 5193
rect 8919 5167 8945 5193
rect 8945 5167 8946 5193
rect 8918 5166 8946 5167
rect 8750 4942 8778 4970
rect 8152 4325 8180 4326
rect 8152 4299 8153 4325
rect 8153 4299 8179 4325
rect 8179 4299 8180 4325
rect 8152 4298 8180 4299
rect 8204 4325 8232 4326
rect 8204 4299 8205 4325
rect 8205 4299 8231 4325
rect 8231 4299 8232 4325
rect 8204 4298 8232 4299
rect 8256 4325 8284 4326
rect 8256 4299 8257 4325
rect 8257 4299 8283 4325
rect 8283 4299 8284 4325
rect 8256 4298 8284 4299
rect 7182 3430 7210 3458
rect 7074 3149 7102 3150
rect 7074 3123 7075 3149
rect 7075 3123 7101 3149
rect 7101 3123 7102 3149
rect 7074 3122 7102 3123
rect 7126 3149 7154 3150
rect 7126 3123 7127 3149
rect 7127 3123 7153 3149
rect 7153 3123 7154 3149
rect 7126 3122 7154 3123
rect 7178 3149 7206 3150
rect 7178 3123 7179 3149
rect 7179 3123 7205 3149
rect 7205 3123 7206 3149
rect 7178 3122 7206 3123
rect 7462 3065 7490 3066
rect 7462 3039 7463 3065
rect 7463 3039 7489 3065
rect 7489 3039 7490 3065
rect 7462 3038 7490 3039
rect 7350 2982 7378 3010
rect 6902 2953 6930 2954
rect 6902 2927 6903 2953
rect 6903 2927 6929 2953
rect 6929 2927 6930 2953
rect 6902 2926 6930 2927
rect 7070 2897 7098 2898
rect 7070 2871 7071 2897
rect 7071 2871 7097 2897
rect 7097 2871 7098 2897
rect 7070 2870 7098 2871
rect 7182 2897 7210 2898
rect 7182 2871 7183 2897
rect 7183 2871 7209 2897
rect 7209 2871 7210 2897
rect 7182 2870 7210 2871
rect 7294 2673 7322 2674
rect 7294 2647 7295 2673
rect 7295 2647 7321 2673
rect 7321 2647 7322 2673
rect 7294 2646 7322 2647
rect 2926 2561 2954 2562
rect 2926 2535 2927 2561
rect 2927 2535 2953 2561
rect 2953 2535 2954 2561
rect 2926 2534 2954 2535
rect 7854 4185 7882 4186
rect 7854 4159 7855 4185
rect 7855 4159 7881 4185
rect 7881 4159 7882 4185
rect 7854 4158 7882 4159
rect 8302 3710 8330 3738
rect 7910 3654 7938 3682
rect 8152 3541 8180 3542
rect 8152 3515 8153 3541
rect 8153 3515 8179 3541
rect 8179 3515 8180 3541
rect 8152 3514 8180 3515
rect 8204 3541 8232 3542
rect 8204 3515 8205 3541
rect 8205 3515 8231 3541
rect 8231 3515 8232 3541
rect 8204 3514 8232 3515
rect 8256 3541 8284 3542
rect 8256 3515 8257 3541
rect 8257 3515 8283 3541
rect 8283 3515 8284 3541
rect 8256 3514 8284 3515
rect 8190 3318 8218 3346
rect 8190 3038 8218 3066
rect 8134 3009 8162 3010
rect 8134 2983 8135 3009
rect 8135 2983 8161 3009
rect 8161 2983 8162 3009
rect 8134 2982 8162 2983
rect 7518 2926 7546 2954
rect 7742 2953 7770 2954
rect 7742 2927 7743 2953
rect 7743 2927 7769 2953
rect 7769 2927 7770 2953
rect 7742 2926 7770 2927
rect 8750 3681 8778 3682
rect 8750 3655 8751 3681
rect 8751 3655 8777 3681
rect 8777 3655 8778 3681
rect 8750 3654 8778 3655
rect 8694 3318 8722 3346
rect 9030 4969 9058 4970
rect 9030 4943 9031 4969
rect 9031 4943 9057 4969
rect 9057 4943 9058 4969
rect 9030 4942 9058 4943
rect 9230 4717 9258 4718
rect 9230 4691 9231 4717
rect 9231 4691 9257 4717
rect 9257 4691 9258 4717
rect 9230 4690 9258 4691
rect 9282 4717 9310 4718
rect 9282 4691 9283 4717
rect 9283 4691 9309 4717
rect 9309 4691 9310 4717
rect 9282 4690 9310 4691
rect 9334 4717 9362 4718
rect 9334 4691 9335 4717
rect 9335 4691 9361 4717
rect 9361 4691 9362 4717
rect 9334 4690 9362 4691
rect 9230 3933 9258 3934
rect 9230 3907 9231 3933
rect 9231 3907 9257 3933
rect 9257 3907 9258 3933
rect 9230 3906 9258 3907
rect 9282 3933 9310 3934
rect 9282 3907 9283 3933
rect 9283 3907 9309 3933
rect 9309 3907 9310 3933
rect 9282 3906 9310 3907
rect 9334 3933 9362 3934
rect 9334 3907 9335 3933
rect 9335 3907 9361 3933
rect 9361 3907 9362 3933
rect 9334 3906 9362 3907
rect 8918 3766 8946 3794
rect 8750 3206 8778 3234
rect 9030 3206 9058 3234
rect 9230 3149 9258 3150
rect 9230 3123 9231 3149
rect 9231 3123 9257 3149
rect 9257 3123 9258 3149
rect 9230 3122 9258 3123
rect 9282 3149 9310 3150
rect 9282 3123 9283 3149
rect 9283 3123 9309 3149
rect 9309 3123 9310 3149
rect 9282 3122 9310 3123
rect 9334 3149 9362 3150
rect 9334 3123 9335 3149
rect 9335 3123 9361 3149
rect 9361 3123 9362 3149
rect 9334 3122 9362 3123
rect 8806 2982 8834 3010
rect 8638 2926 8666 2954
rect 7406 2814 7434 2842
rect 8918 2814 8946 2842
rect 8152 2757 8180 2758
rect 8152 2731 8153 2757
rect 8153 2731 8179 2757
rect 8179 2731 8180 2757
rect 8152 2730 8180 2731
rect 8204 2757 8232 2758
rect 8204 2731 8205 2757
rect 8205 2731 8231 2757
rect 8231 2731 8232 2757
rect 8204 2730 8232 2731
rect 8256 2757 8284 2758
rect 8256 2731 8257 2757
rect 8257 2731 8283 2757
rect 8283 2731 8284 2757
rect 8256 2730 8284 2731
rect 2762 2365 2790 2366
rect 2762 2339 2763 2365
rect 2763 2339 2789 2365
rect 2789 2339 2790 2365
rect 2762 2338 2790 2339
rect 2814 2365 2842 2366
rect 2814 2339 2815 2365
rect 2815 2339 2841 2365
rect 2841 2339 2842 2365
rect 2814 2338 2842 2339
rect 2866 2365 2894 2366
rect 2866 2339 2867 2365
rect 2867 2339 2893 2365
rect 2893 2339 2894 2365
rect 2866 2338 2894 2339
rect 4918 2365 4946 2366
rect 4918 2339 4919 2365
rect 4919 2339 4945 2365
rect 4945 2339 4946 2365
rect 4918 2338 4946 2339
rect 4970 2365 4998 2366
rect 4970 2339 4971 2365
rect 4971 2339 4997 2365
rect 4997 2339 4998 2365
rect 4970 2338 4998 2339
rect 5022 2365 5050 2366
rect 5022 2339 5023 2365
rect 5023 2339 5049 2365
rect 5049 2339 5050 2365
rect 5022 2338 5050 2339
rect 7074 2365 7102 2366
rect 7074 2339 7075 2365
rect 7075 2339 7101 2365
rect 7101 2339 7102 2365
rect 7074 2338 7102 2339
rect 7126 2365 7154 2366
rect 7126 2339 7127 2365
rect 7127 2339 7153 2365
rect 7153 2339 7154 2365
rect 7126 2338 7154 2339
rect 7178 2365 7206 2366
rect 7178 2339 7179 2365
rect 7179 2339 7205 2365
rect 7205 2339 7206 2365
rect 7178 2338 7206 2339
rect 3840 1973 3868 1974
rect 3840 1947 3841 1973
rect 3841 1947 3867 1973
rect 3867 1947 3868 1973
rect 3840 1946 3868 1947
rect 3892 1973 3920 1974
rect 3892 1947 3893 1973
rect 3893 1947 3919 1973
rect 3919 1947 3920 1973
rect 3892 1946 3920 1947
rect 3944 1973 3972 1974
rect 3944 1947 3945 1973
rect 3945 1947 3971 1973
rect 3971 1947 3972 1973
rect 3944 1946 3972 1947
rect 5996 1973 6024 1974
rect 5996 1947 5997 1973
rect 5997 1947 6023 1973
rect 6023 1947 6024 1973
rect 5996 1946 6024 1947
rect 6048 1973 6076 1974
rect 6048 1947 6049 1973
rect 6049 1947 6075 1973
rect 6075 1947 6076 1973
rect 6048 1946 6076 1947
rect 6100 1973 6128 1974
rect 6100 1947 6101 1973
rect 6101 1947 6127 1973
rect 6127 1947 6128 1973
rect 6100 1946 6128 1947
rect 8152 1973 8180 1974
rect 8152 1947 8153 1973
rect 8153 1947 8179 1973
rect 8179 1947 8180 1973
rect 8152 1946 8180 1947
rect 8204 1973 8232 1974
rect 8204 1947 8205 1973
rect 8205 1947 8231 1973
rect 8231 1947 8232 1973
rect 8204 1946 8232 1947
rect 8256 1973 8284 1974
rect 8256 1947 8257 1973
rect 8257 1947 8283 1973
rect 8283 1947 8284 1973
rect 8256 1946 8284 1947
rect 9230 2365 9258 2366
rect 9230 2339 9231 2365
rect 9231 2339 9257 2365
rect 9257 2339 9258 2365
rect 9230 2338 9258 2339
rect 9282 2365 9310 2366
rect 9282 2339 9283 2365
rect 9283 2339 9309 2365
rect 9309 2339 9310 2365
rect 9282 2338 9310 2339
rect 9334 2365 9362 2366
rect 9334 2339 9335 2365
rect 9335 2339 9361 2365
rect 9361 2339 9362 2365
rect 9334 2338 9362 2339
rect 8806 1638 8834 1666
rect 9086 1638 9114 1666
rect 2762 1581 2790 1582
rect 2762 1555 2763 1581
rect 2763 1555 2789 1581
rect 2789 1555 2790 1581
rect 2762 1554 2790 1555
rect 2814 1581 2842 1582
rect 2814 1555 2815 1581
rect 2815 1555 2841 1581
rect 2841 1555 2842 1581
rect 2814 1554 2842 1555
rect 2866 1581 2894 1582
rect 2866 1555 2867 1581
rect 2867 1555 2893 1581
rect 2893 1555 2894 1581
rect 2866 1554 2894 1555
rect 4918 1581 4946 1582
rect 4918 1555 4919 1581
rect 4919 1555 4945 1581
rect 4945 1555 4946 1581
rect 4918 1554 4946 1555
rect 4970 1581 4998 1582
rect 4970 1555 4971 1581
rect 4971 1555 4997 1581
rect 4997 1555 4998 1581
rect 4970 1554 4998 1555
rect 5022 1581 5050 1582
rect 5022 1555 5023 1581
rect 5023 1555 5049 1581
rect 5049 1555 5050 1581
rect 5022 1554 5050 1555
rect 7074 1581 7102 1582
rect 7074 1555 7075 1581
rect 7075 1555 7101 1581
rect 7101 1555 7102 1581
rect 7074 1554 7102 1555
rect 7126 1581 7154 1582
rect 7126 1555 7127 1581
rect 7127 1555 7153 1581
rect 7153 1555 7154 1581
rect 7126 1554 7154 1555
rect 7178 1581 7206 1582
rect 7178 1555 7179 1581
rect 7179 1555 7205 1581
rect 7205 1555 7206 1581
rect 7178 1554 7206 1555
rect 9230 1581 9258 1582
rect 9230 1555 9231 1581
rect 9231 1555 9257 1581
rect 9257 1555 9258 1581
rect 9230 1554 9258 1555
rect 9282 1581 9310 1582
rect 9282 1555 9283 1581
rect 9283 1555 9309 1581
rect 9309 1555 9310 1581
rect 9282 1554 9310 1555
rect 9334 1581 9362 1582
rect 9334 1555 9335 1581
rect 9335 1555 9361 1581
rect 9361 1555 9362 1581
rect 9334 1554 9362 1555
rect 9086 1246 9114 1274
rect 966 630 994 658
<< metal3 >>
rect 0 9226 400 9240
rect 0 9198 1190 9226
rect 1218 9198 1223 9226
rect 0 9184 400 9198
rect 9600 8666 10000 8680
rect 7457 8638 7462 8666
rect 7490 8638 10000 8666
rect 9600 8624 10000 8638
rect 1679 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1821 8246
rect 3835 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3977 8246
rect 5991 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6133 8246
rect 8147 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8289 8246
rect 7401 8022 7406 8050
rect 7434 8022 8358 8050
rect 8386 8022 8582 8050
rect 8610 8022 8615 8050
rect 0 7994 400 8008
rect 0 7966 854 7994
rect 882 7966 1582 7994
rect 1610 7966 1615 7994
rect 0 7952 400 7966
rect 2757 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2899 7854
rect 4913 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5055 7854
rect 7069 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7211 7854
rect 9225 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9367 7854
rect 1073 7742 1078 7770
rect 1106 7742 1190 7770
rect 1218 7742 1223 7770
rect 1465 7630 1470 7658
rect 1498 7630 3150 7658
rect 3178 7630 3183 7658
rect 2865 7574 2870 7602
rect 2898 7574 4102 7602
rect 4130 7574 4135 7602
rect 2473 7518 2478 7546
rect 2506 7518 4438 7546
rect 4466 7518 4471 7546
rect 1679 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1821 7462
rect 3835 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3977 7462
rect 5991 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6133 7462
rect 8147 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8289 7462
rect 2977 7294 2982 7322
rect 3010 7294 3598 7322
rect 3626 7294 3631 7322
rect 3761 7294 3766 7322
rect 3794 7294 4270 7322
rect 4298 7294 6174 7322
rect 6202 7294 6207 7322
rect 3257 7238 3262 7266
rect 3290 7238 3654 7266
rect 3682 7238 3687 7266
rect 4186 7238 6958 7266
rect 6986 7238 7518 7266
rect 7546 7238 7551 7266
rect 4186 7210 4214 7238
rect 3313 7182 3318 7210
rect 3346 7182 4214 7210
rect 4489 7182 4494 7210
rect 4522 7182 5110 7210
rect 5138 7182 5143 7210
rect 4937 7126 4942 7154
rect 4970 7126 5866 7154
rect 5838 7098 5866 7126
rect 5833 7070 5838 7098
rect 5866 7070 6510 7098
rect 6538 7070 6543 7098
rect 2757 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2899 7070
rect 4913 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5055 7070
rect 7069 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7211 7070
rect 9225 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9367 7070
rect 2641 6958 2646 6986
rect 2674 6958 3206 6986
rect 3234 6958 3542 6986
rect 3570 6958 3878 6986
rect 3906 6958 8470 6986
rect 8498 6958 8503 6986
rect 5609 6902 5614 6930
rect 5642 6902 7630 6930
rect 7658 6902 7663 6930
rect 5161 6846 5166 6874
rect 5194 6846 6118 6874
rect 6146 6846 6151 6874
rect 3985 6790 3990 6818
rect 4018 6790 4158 6818
rect 4186 6790 5334 6818
rect 5362 6790 5367 6818
rect 0 6762 400 6776
rect 0 6734 854 6762
rect 882 6734 1246 6762
rect 1274 6734 1279 6762
rect 5889 6734 5894 6762
rect 5922 6734 7546 6762
rect 0 6720 400 6734
rect 7518 6706 7546 6734
rect 7518 6678 7686 6706
rect 7714 6678 7719 6706
rect 1679 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1821 6678
rect 3835 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3977 6678
rect 5991 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6133 6678
rect 8147 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8289 6678
rect 6169 6566 6174 6594
rect 6202 6566 6790 6594
rect 6818 6566 6823 6594
rect 4186 6510 7574 6538
rect 7602 6510 7607 6538
rect 4186 6482 4214 6510
rect 3649 6454 3654 6482
rect 3682 6454 4214 6482
rect 7457 6454 7462 6482
rect 7490 6454 7966 6482
rect 7994 6454 7999 6482
rect 4186 6398 5054 6426
rect 5082 6398 5087 6426
rect 2757 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2899 6286
rect 4186 6202 4214 6398
rect 4657 6342 4662 6370
rect 4690 6342 6342 6370
rect 6370 6342 6622 6370
rect 6650 6342 6655 6370
rect 6841 6342 6846 6370
rect 6874 6342 7238 6370
rect 7266 6342 7271 6370
rect 5945 6286 5950 6314
rect 5978 6286 6902 6314
rect 6930 6286 6935 6314
rect 4913 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5055 6286
rect 7069 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7211 6286
rect 9225 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9367 6286
rect 5502 6230 6202 6258
rect 5502 6202 5530 6230
rect 6174 6202 6202 6230
rect 9600 6202 10000 6216
rect 1073 6174 1078 6202
rect 1106 6174 1974 6202
rect 2002 6174 2478 6202
rect 2506 6174 2511 6202
rect 3481 6174 3486 6202
rect 3514 6174 4214 6202
rect 4242 6174 4247 6202
rect 4489 6174 4494 6202
rect 4522 6174 4830 6202
rect 4858 6174 5530 6202
rect 5609 6174 5614 6202
rect 5642 6174 5838 6202
rect 5866 6174 5871 6202
rect 6174 6174 7014 6202
rect 7042 6174 7238 6202
rect 7266 6174 7271 6202
rect 8969 6174 8974 6202
rect 9002 6174 10000 6202
rect 9600 6160 10000 6174
rect 4545 6118 4550 6146
rect 4578 6118 4886 6146
rect 4914 6118 5222 6146
rect 5250 6118 5255 6146
rect 6001 6118 6006 6146
rect 6034 6118 6734 6146
rect 6762 6118 6767 6146
rect 1577 6062 1582 6090
rect 1610 6062 2982 6090
rect 3010 6062 3318 6090
rect 3346 6062 3351 6090
rect 4377 6062 4382 6090
rect 4410 6062 4942 6090
rect 4970 6062 6062 6090
rect 6090 6062 6095 6090
rect 6225 6062 6230 6090
rect 6258 6062 6846 6090
rect 6874 6062 6879 6090
rect 6953 6062 6958 6090
rect 6986 6062 7406 6090
rect 7434 6062 7910 6090
rect 7938 6062 7943 6090
rect 5105 6006 5110 6034
rect 5138 6006 5670 6034
rect 5698 6006 5703 6034
rect 6673 5950 6678 5978
rect 6706 5950 7574 5978
rect 7602 5950 7607 5978
rect 7737 5950 7742 5978
rect 7770 5950 7966 5978
rect 7994 5950 7999 5978
rect 2361 5894 2366 5922
rect 2394 5894 2534 5922
rect 2562 5894 3318 5922
rect 3346 5894 3351 5922
rect 5329 5894 5334 5922
rect 5362 5894 5894 5922
rect 5922 5894 5927 5922
rect 6790 5894 7686 5922
rect 7714 5894 7719 5922
rect 1679 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1821 5894
rect 3835 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3977 5894
rect 5991 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6133 5894
rect 6790 5810 6818 5894
rect 8147 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8289 5894
rect 6785 5782 6790 5810
rect 6818 5782 6823 5810
rect 6561 5726 6566 5754
rect 6594 5726 7574 5754
rect 7602 5726 7607 5754
rect 8073 5726 8078 5754
rect 8106 5726 9086 5754
rect 9114 5726 9119 5754
rect 6617 5670 6622 5698
rect 6650 5670 6846 5698
rect 6874 5670 6879 5698
rect 6393 5614 6398 5642
rect 6426 5614 7126 5642
rect 7154 5614 7159 5642
rect 7457 5614 7462 5642
rect 7490 5614 8022 5642
rect 8050 5614 8055 5642
rect 1185 5558 1190 5586
rect 1218 5558 2142 5586
rect 2170 5558 2175 5586
rect 4545 5558 4550 5586
rect 4578 5558 5222 5586
rect 5250 5558 5255 5586
rect 6958 5558 7182 5586
rect 7210 5558 7215 5586
rect 0 5530 400 5544
rect 6958 5530 6986 5558
rect 0 5502 854 5530
rect 882 5502 1246 5530
rect 1274 5502 1279 5530
rect 6953 5502 6958 5530
rect 6986 5502 6991 5530
rect 0 5488 400 5502
rect 2757 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2899 5502
rect 4913 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5055 5502
rect 7069 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7211 5502
rect 9225 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9367 5502
rect 1129 5390 1134 5418
rect 1162 5390 2814 5418
rect 2842 5390 3430 5418
rect 3458 5390 4102 5418
rect 4130 5390 4135 5418
rect 4489 5390 4494 5418
rect 4522 5390 5166 5418
rect 5194 5390 5199 5418
rect 2305 5334 2310 5362
rect 2338 5334 2646 5362
rect 2674 5334 2679 5362
rect 5833 5334 5838 5362
rect 5866 5334 6174 5362
rect 6202 5334 6207 5362
rect 7009 5278 7014 5306
rect 7042 5278 8078 5306
rect 8106 5278 8111 5306
rect 1017 5222 1022 5250
rect 1050 5222 1414 5250
rect 1442 5222 1447 5250
rect 4825 5222 4830 5250
rect 4858 5222 6342 5250
rect 6370 5222 6375 5250
rect 2193 5166 2198 5194
rect 2226 5166 2590 5194
rect 2618 5166 4718 5194
rect 4746 5166 4751 5194
rect 7345 5166 7350 5194
rect 7378 5166 8918 5194
rect 8946 5166 8951 5194
rect 3201 5110 3206 5138
rect 3234 5110 3374 5138
rect 3402 5110 3407 5138
rect 1679 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1821 5110
rect 3835 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3977 5110
rect 5991 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6133 5110
rect 8147 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8289 5110
rect 1862 5054 2478 5082
rect 2506 5054 2511 5082
rect 2641 5054 2646 5082
rect 2674 5054 3150 5082
rect 3178 5054 3183 5082
rect 1862 5026 1890 5054
rect 1633 4998 1638 5026
rect 1666 4998 1890 5026
rect 6449 4998 6454 5026
rect 6482 4998 7014 5026
rect 7042 4998 7047 5026
rect 7121 4998 7126 5026
rect 7154 4998 7686 5026
rect 7714 4998 8022 5026
rect 8050 4998 8055 5026
rect 1465 4942 1470 4970
rect 1498 4942 1694 4970
rect 1722 4942 1727 4970
rect 3257 4942 3262 4970
rect 3290 4942 3542 4970
rect 3570 4942 3575 4970
rect 4321 4942 4326 4970
rect 4354 4942 6510 4970
rect 6538 4942 6734 4970
rect 6762 4942 6767 4970
rect 7233 4942 7238 4970
rect 7266 4942 7742 4970
rect 7770 4942 8302 4970
rect 8330 4942 8335 4970
rect 8745 4942 8750 4970
rect 8778 4942 9030 4970
rect 9058 4942 9063 4970
rect 2529 4886 2534 4914
rect 2562 4886 4214 4914
rect 4825 4886 4830 4914
rect 4858 4886 5446 4914
rect 5474 4886 5479 4914
rect 4186 4858 4214 4886
rect 2025 4830 2030 4858
rect 2058 4830 2422 4858
rect 2450 4830 2926 4858
rect 2954 4830 2959 4858
rect 4186 4830 4774 4858
rect 4802 4830 4807 4858
rect 4886 4802 4914 4886
rect 8750 4858 8778 4942
rect 5273 4830 5278 4858
rect 5306 4830 8778 4858
rect 4041 4774 4046 4802
rect 4074 4774 4382 4802
rect 4410 4774 4415 4802
rect 4489 4774 4494 4802
rect 4522 4774 4914 4802
rect 6673 4774 6678 4802
rect 6706 4774 6902 4802
rect 6930 4774 6935 4802
rect 4433 4718 4438 4746
rect 4466 4718 4830 4746
rect 4858 4718 4863 4746
rect 2757 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2899 4718
rect 4913 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5055 4718
rect 7069 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7211 4718
rect 9225 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9367 4718
rect 3313 4606 3318 4634
rect 3346 4606 5502 4634
rect 5530 4606 5535 4634
rect 6841 4606 6846 4634
rect 6874 4606 7462 4634
rect 7490 4606 7495 4634
rect 1409 4550 1414 4578
rect 1442 4550 2366 4578
rect 2394 4550 2399 4578
rect 4545 4550 4550 4578
rect 4578 4550 5894 4578
rect 5922 4550 6174 4578
rect 6202 4550 6207 4578
rect 1521 4494 1526 4522
rect 1554 4494 2142 4522
rect 2170 4494 2175 4522
rect 2529 4494 2534 4522
rect 2562 4494 3318 4522
rect 3346 4494 4326 4522
rect 4354 4494 4359 4522
rect 4489 4494 4494 4522
rect 4522 4494 4830 4522
rect 4858 4494 4863 4522
rect 4494 4466 4522 4494
rect 4209 4438 4214 4466
rect 4242 4438 4522 4466
rect 1465 4382 1470 4410
rect 1498 4382 2086 4410
rect 2114 4382 2119 4410
rect 2305 4382 2310 4410
rect 2338 4382 3206 4410
rect 3234 4382 3239 4410
rect 0 4298 400 4312
rect 1679 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1821 4326
rect 3835 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3977 4326
rect 5991 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6133 4326
rect 8147 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8289 4326
rect 0 4270 854 4298
rect 882 4270 1246 4298
rect 1274 4270 1279 4298
rect 5049 4270 5054 4298
rect 5082 4270 5726 4298
rect 5754 4270 5759 4298
rect 0 4256 400 4270
rect 3817 4214 3822 4242
rect 3850 4214 5334 4242
rect 5362 4214 5367 4242
rect 4265 4158 4270 4186
rect 4298 4158 4886 4186
rect 4914 4158 5222 4186
rect 5250 4158 5255 4186
rect 5665 4158 5670 4186
rect 5698 4158 5894 4186
rect 5922 4158 6622 4186
rect 6650 4158 6655 4186
rect 7401 4158 7406 4186
rect 7434 4158 7854 4186
rect 7882 4158 7887 4186
rect 6230 4130 6258 4158
rect 5105 4102 5110 4130
rect 5138 4102 5558 4130
rect 5586 4102 5591 4130
rect 6225 4102 6230 4130
rect 6258 4102 6263 4130
rect 6449 4102 6454 4130
rect 6482 4102 6790 4130
rect 6818 4102 6823 4130
rect 5329 4046 5334 4074
rect 5362 4046 5894 4074
rect 5922 4046 5927 4074
rect 2921 3990 2926 4018
rect 2954 3990 4158 4018
rect 4186 3990 4191 4018
rect 6902 3990 7238 4018
rect 7266 3990 7271 4018
rect 6902 3962 6930 3990
rect 6785 3934 6790 3962
rect 6818 3934 6930 3962
rect 2757 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2899 3934
rect 4913 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5055 3934
rect 7069 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7211 3934
rect 9225 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9367 3934
rect 2697 3822 2702 3850
rect 2730 3822 3374 3850
rect 3402 3822 3407 3850
rect 4489 3822 4494 3850
rect 4522 3822 5110 3850
rect 5138 3822 5143 3850
rect 6169 3822 6174 3850
rect 6202 3822 6734 3850
rect 6762 3822 7070 3850
rect 7098 3822 7103 3850
rect 3201 3766 3206 3794
rect 3234 3766 4718 3794
rect 4746 3766 4751 3794
rect 5553 3766 5558 3794
rect 5586 3766 8918 3794
rect 8946 3766 8951 3794
rect 7014 3738 7042 3766
rect 9600 3738 10000 3752
rect 2977 3710 2982 3738
rect 3010 3710 3318 3738
rect 3346 3710 3351 3738
rect 3873 3710 3878 3738
rect 3906 3710 4886 3738
rect 4914 3710 4919 3738
rect 6953 3710 6958 3738
rect 6986 3710 7042 3738
rect 8297 3710 8302 3738
rect 8330 3710 10000 3738
rect 9600 3696 10000 3710
rect 7905 3654 7910 3682
rect 7938 3654 8750 3682
rect 8778 3654 8783 3682
rect 2865 3598 2870 3626
rect 2898 3598 3430 3626
rect 3458 3598 3463 3626
rect 3761 3598 3766 3626
rect 3794 3598 4270 3626
rect 4298 3598 4830 3626
rect 4858 3598 5838 3626
rect 5866 3598 7014 3626
rect 7042 3598 7047 3626
rect 1679 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1821 3542
rect 3835 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3977 3542
rect 5991 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6133 3542
rect 8147 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8289 3542
rect 6225 3430 6230 3458
rect 6258 3430 7182 3458
rect 7210 3430 7215 3458
rect 6281 3374 6286 3402
rect 6314 3374 6762 3402
rect 1465 3318 1470 3346
rect 1498 3318 3038 3346
rect 3066 3318 3071 3346
rect 4993 3318 4998 3346
rect 5026 3318 6174 3346
rect 6202 3318 6207 3346
rect 6734 3290 6762 3374
rect 8185 3318 8190 3346
rect 8218 3318 8694 3346
rect 8722 3318 8727 3346
rect 5217 3262 5222 3290
rect 5250 3262 6398 3290
rect 6426 3262 6431 3290
rect 6729 3262 6734 3290
rect 6762 3262 6767 3290
rect 6841 3206 6846 3234
rect 6874 3206 8750 3234
rect 8778 3206 9030 3234
rect 9058 3206 9063 3234
rect 2757 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2899 3150
rect 4913 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5055 3150
rect 7069 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7211 3150
rect 9225 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9367 3150
rect 0 3066 400 3080
rect 0 3038 854 3066
rect 882 3038 1246 3066
rect 1274 3038 1279 3066
rect 7457 3038 7462 3066
rect 7490 3038 8190 3066
rect 8218 3038 8223 3066
rect 0 3024 400 3038
rect 7345 2982 7350 3010
rect 7378 2982 8134 3010
rect 8162 2982 8806 3010
rect 8834 2982 8839 3010
rect 6897 2926 6902 2954
rect 6930 2926 7518 2954
rect 7546 2926 7551 2954
rect 7737 2926 7742 2954
rect 7770 2926 8638 2954
rect 8666 2926 8671 2954
rect 7742 2898 7770 2926
rect 5777 2870 5782 2898
rect 5810 2870 7070 2898
rect 7098 2870 7103 2898
rect 7177 2870 7182 2898
rect 7210 2870 7770 2898
rect 6393 2814 6398 2842
rect 6426 2814 7406 2842
rect 7434 2814 8918 2842
rect 8946 2814 8951 2842
rect 1679 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1821 2758
rect 3835 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3977 2758
rect 5991 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6133 2758
rect 8147 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8289 2758
rect 6169 2646 6174 2674
rect 6202 2646 7294 2674
rect 7322 2646 7327 2674
rect 1017 2534 1022 2562
rect 1050 2534 2926 2562
rect 2954 2534 2959 2562
rect 2757 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2899 2366
rect 4913 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5055 2366
rect 7069 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7211 2366
rect 9225 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9367 2366
rect 849 2086 854 2114
rect 882 2086 1246 2114
rect 1274 2086 1279 2114
rect 1679 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1821 1974
rect 3835 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3977 1974
rect 5991 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6133 1974
rect 8147 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8289 1974
rect 0 1834 400 1848
rect 0 1806 854 1834
rect 882 1806 887 1834
rect 0 1792 400 1806
rect 8801 1638 8806 1666
rect 8834 1638 9086 1666
rect 9114 1638 9119 1666
rect 2757 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2899 1582
rect 4913 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5055 1582
rect 7069 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7211 1582
rect 9225 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9367 1582
rect 9600 1274 10000 1288
rect 9081 1246 9086 1274
rect 9114 1246 10000 1274
rect 9600 1232 10000 1246
rect 462 630 966 658
rect 994 630 999 658
rect 0 602 400 616
rect 462 602 490 630
rect 0 574 490 602
rect 0 560 400 574
<< via3 >>
rect 1684 8218 1712 8246
rect 1736 8218 1764 8246
rect 1788 8218 1816 8246
rect 3840 8218 3868 8246
rect 3892 8218 3920 8246
rect 3944 8218 3972 8246
rect 5996 8218 6024 8246
rect 6048 8218 6076 8246
rect 6100 8218 6128 8246
rect 8152 8218 8180 8246
rect 8204 8218 8232 8246
rect 8256 8218 8284 8246
rect 2762 7826 2790 7854
rect 2814 7826 2842 7854
rect 2866 7826 2894 7854
rect 4918 7826 4946 7854
rect 4970 7826 4998 7854
rect 5022 7826 5050 7854
rect 7074 7826 7102 7854
rect 7126 7826 7154 7854
rect 7178 7826 7206 7854
rect 9230 7826 9258 7854
rect 9282 7826 9310 7854
rect 9334 7826 9362 7854
rect 1684 7434 1712 7462
rect 1736 7434 1764 7462
rect 1788 7434 1816 7462
rect 3840 7434 3868 7462
rect 3892 7434 3920 7462
rect 3944 7434 3972 7462
rect 5996 7434 6024 7462
rect 6048 7434 6076 7462
rect 6100 7434 6128 7462
rect 8152 7434 8180 7462
rect 8204 7434 8232 7462
rect 8256 7434 8284 7462
rect 2762 7042 2790 7070
rect 2814 7042 2842 7070
rect 2866 7042 2894 7070
rect 4918 7042 4946 7070
rect 4970 7042 4998 7070
rect 5022 7042 5050 7070
rect 7074 7042 7102 7070
rect 7126 7042 7154 7070
rect 7178 7042 7206 7070
rect 9230 7042 9258 7070
rect 9282 7042 9310 7070
rect 9334 7042 9362 7070
rect 1684 6650 1712 6678
rect 1736 6650 1764 6678
rect 1788 6650 1816 6678
rect 3840 6650 3868 6678
rect 3892 6650 3920 6678
rect 3944 6650 3972 6678
rect 5996 6650 6024 6678
rect 6048 6650 6076 6678
rect 6100 6650 6128 6678
rect 8152 6650 8180 6678
rect 8204 6650 8232 6678
rect 8256 6650 8284 6678
rect 2762 6258 2790 6286
rect 2814 6258 2842 6286
rect 2866 6258 2894 6286
rect 4918 6258 4946 6286
rect 4970 6258 4998 6286
rect 5022 6258 5050 6286
rect 7074 6258 7102 6286
rect 7126 6258 7154 6286
rect 7178 6258 7206 6286
rect 9230 6258 9258 6286
rect 9282 6258 9310 6286
rect 9334 6258 9362 6286
rect 1684 5866 1712 5894
rect 1736 5866 1764 5894
rect 1788 5866 1816 5894
rect 3840 5866 3868 5894
rect 3892 5866 3920 5894
rect 3944 5866 3972 5894
rect 5996 5866 6024 5894
rect 6048 5866 6076 5894
rect 6100 5866 6128 5894
rect 8152 5866 8180 5894
rect 8204 5866 8232 5894
rect 8256 5866 8284 5894
rect 2762 5474 2790 5502
rect 2814 5474 2842 5502
rect 2866 5474 2894 5502
rect 4918 5474 4946 5502
rect 4970 5474 4998 5502
rect 5022 5474 5050 5502
rect 7074 5474 7102 5502
rect 7126 5474 7154 5502
rect 7178 5474 7206 5502
rect 9230 5474 9258 5502
rect 9282 5474 9310 5502
rect 9334 5474 9362 5502
rect 1684 5082 1712 5110
rect 1736 5082 1764 5110
rect 1788 5082 1816 5110
rect 3840 5082 3868 5110
rect 3892 5082 3920 5110
rect 3944 5082 3972 5110
rect 5996 5082 6024 5110
rect 6048 5082 6076 5110
rect 6100 5082 6128 5110
rect 8152 5082 8180 5110
rect 8204 5082 8232 5110
rect 8256 5082 8284 5110
rect 2762 4690 2790 4718
rect 2814 4690 2842 4718
rect 2866 4690 2894 4718
rect 4918 4690 4946 4718
rect 4970 4690 4998 4718
rect 5022 4690 5050 4718
rect 7074 4690 7102 4718
rect 7126 4690 7154 4718
rect 7178 4690 7206 4718
rect 9230 4690 9258 4718
rect 9282 4690 9310 4718
rect 9334 4690 9362 4718
rect 1684 4298 1712 4326
rect 1736 4298 1764 4326
rect 1788 4298 1816 4326
rect 3840 4298 3868 4326
rect 3892 4298 3920 4326
rect 3944 4298 3972 4326
rect 5996 4298 6024 4326
rect 6048 4298 6076 4326
rect 6100 4298 6128 4326
rect 8152 4298 8180 4326
rect 8204 4298 8232 4326
rect 8256 4298 8284 4326
rect 2762 3906 2790 3934
rect 2814 3906 2842 3934
rect 2866 3906 2894 3934
rect 4918 3906 4946 3934
rect 4970 3906 4998 3934
rect 5022 3906 5050 3934
rect 7074 3906 7102 3934
rect 7126 3906 7154 3934
rect 7178 3906 7206 3934
rect 9230 3906 9258 3934
rect 9282 3906 9310 3934
rect 9334 3906 9362 3934
rect 1684 3514 1712 3542
rect 1736 3514 1764 3542
rect 1788 3514 1816 3542
rect 3840 3514 3868 3542
rect 3892 3514 3920 3542
rect 3944 3514 3972 3542
rect 5996 3514 6024 3542
rect 6048 3514 6076 3542
rect 6100 3514 6128 3542
rect 8152 3514 8180 3542
rect 8204 3514 8232 3542
rect 8256 3514 8284 3542
rect 2762 3122 2790 3150
rect 2814 3122 2842 3150
rect 2866 3122 2894 3150
rect 4918 3122 4946 3150
rect 4970 3122 4998 3150
rect 5022 3122 5050 3150
rect 7074 3122 7102 3150
rect 7126 3122 7154 3150
rect 7178 3122 7206 3150
rect 9230 3122 9258 3150
rect 9282 3122 9310 3150
rect 9334 3122 9362 3150
rect 1684 2730 1712 2758
rect 1736 2730 1764 2758
rect 1788 2730 1816 2758
rect 3840 2730 3868 2758
rect 3892 2730 3920 2758
rect 3944 2730 3972 2758
rect 5996 2730 6024 2758
rect 6048 2730 6076 2758
rect 6100 2730 6128 2758
rect 8152 2730 8180 2758
rect 8204 2730 8232 2758
rect 8256 2730 8284 2758
rect 2762 2338 2790 2366
rect 2814 2338 2842 2366
rect 2866 2338 2894 2366
rect 4918 2338 4946 2366
rect 4970 2338 4998 2366
rect 5022 2338 5050 2366
rect 7074 2338 7102 2366
rect 7126 2338 7154 2366
rect 7178 2338 7206 2366
rect 9230 2338 9258 2366
rect 9282 2338 9310 2366
rect 9334 2338 9362 2366
rect 1684 1946 1712 1974
rect 1736 1946 1764 1974
rect 1788 1946 1816 1974
rect 3840 1946 3868 1974
rect 3892 1946 3920 1974
rect 3944 1946 3972 1974
rect 5996 1946 6024 1974
rect 6048 1946 6076 1974
rect 6100 1946 6128 1974
rect 8152 1946 8180 1974
rect 8204 1946 8232 1974
rect 8256 1946 8284 1974
rect 2762 1554 2790 1582
rect 2814 1554 2842 1582
rect 2866 1554 2894 1582
rect 4918 1554 4946 1582
rect 4970 1554 4998 1582
rect 5022 1554 5050 1582
rect 7074 1554 7102 1582
rect 7126 1554 7154 1582
rect 7178 1554 7206 1582
rect 9230 1554 9258 1582
rect 9282 1554 9310 1582
rect 9334 1554 9362 1582
<< metal4 >>
rect 1670 8246 1830 8262
rect 1670 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1830 8246
rect 1670 7462 1830 8218
rect 1670 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1830 7462
rect 1670 6678 1830 7434
rect 1670 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1830 6678
rect 1670 5894 1830 6650
rect 1670 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1830 5894
rect 1670 5110 1830 5866
rect 1670 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1830 5110
rect 1670 4326 1830 5082
rect 1670 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1830 4326
rect 1670 3542 1830 4298
rect 1670 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1830 3542
rect 1670 2758 1830 3514
rect 1670 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1830 2758
rect 1670 1974 1830 2730
rect 1670 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1830 1974
rect 1670 1538 1830 1946
rect 2748 7854 2908 8262
rect 2748 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2908 7854
rect 2748 7070 2908 7826
rect 2748 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2908 7070
rect 2748 6286 2908 7042
rect 2748 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2908 6286
rect 2748 5502 2908 6258
rect 2748 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2908 5502
rect 2748 4718 2908 5474
rect 2748 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2908 4718
rect 2748 3934 2908 4690
rect 2748 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2908 3934
rect 2748 3150 2908 3906
rect 2748 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2908 3150
rect 2748 2366 2908 3122
rect 2748 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2908 2366
rect 2748 1582 2908 2338
rect 2748 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2908 1582
rect 2748 1538 2908 1554
rect 3826 8246 3986 8262
rect 3826 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3986 8246
rect 3826 7462 3986 8218
rect 3826 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3986 7462
rect 3826 6678 3986 7434
rect 3826 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3986 6678
rect 3826 5894 3986 6650
rect 3826 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3986 5894
rect 3826 5110 3986 5866
rect 3826 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3986 5110
rect 3826 4326 3986 5082
rect 3826 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3986 4326
rect 3826 3542 3986 4298
rect 3826 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3986 3542
rect 3826 2758 3986 3514
rect 3826 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3986 2758
rect 3826 1974 3986 2730
rect 3826 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3986 1974
rect 3826 1538 3986 1946
rect 4904 7854 5064 8262
rect 4904 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5064 7854
rect 4904 7070 5064 7826
rect 4904 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5064 7070
rect 4904 6286 5064 7042
rect 4904 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5064 6286
rect 4904 5502 5064 6258
rect 4904 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5064 5502
rect 4904 4718 5064 5474
rect 4904 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5064 4718
rect 4904 3934 5064 4690
rect 4904 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5064 3934
rect 4904 3150 5064 3906
rect 4904 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5064 3150
rect 4904 2366 5064 3122
rect 4904 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5064 2366
rect 4904 1582 5064 2338
rect 4904 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5064 1582
rect 4904 1538 5064 1554
rect 5982 8246 6142 8262
rect 5982 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6142 8246
rect 5982 7462 6142 8218
rect 5982 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6142 7462
rect 5982 6678 6142 7434
rect 5982 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6142 6678
rect 5982 5894 6142 6650
rect 5982 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6142 5894
rect 5982 5110 6142 5866
rect 5982 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6142 5110
rect 5982 4326 6142 5082
rect 5982 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6142 4326
rect 5982 3542 6142 4298
rect 5982 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6142 3542
rect 5982 2758 6142 3514
rect 5982 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6142 2758
rect 5982 1974 6142 2730
rect 5982 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6142 1974
rect 5982 1538 6142 1946
rect 7060 7854 7220 8262
rect 7060 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7220 7854
rect 7060 7070 7220 7826
rect 7060 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7220 7070
rect 7060 6286 7220 7042
rect 7060 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7220 6286
rect 7060 5502 7220 6258
rect 7060 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7220 5502
rect 7060 4718 7220 5474
rect 7060 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7220 4718
rect 7060 3934 7220 4690
rect 7060 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7220 3934
rect 7060 3150 7220 3906
rect 7060 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7220 3150
rect 7060 2366 7220 3122
rect 7060 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7220 2366
rect 7060 1582 7220 2338
rect 7060 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7220 1582
rect 7060 1538 7220 1554
rect 8138 8246 8298 8262
rect 8138 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8298 8246
rect 8138 7462 8298 8218
rect 8138 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8298 7462
rect 8138 6678 8298 7434
rect 8138 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8298 6678
rect 8138 5894 8298 6650
rect 8138 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8298 5894
rect 8138 5110 8298 5866
rect 8138 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8298 5110
rect 8138 4326 8298 5082
rect 8138 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8298 4326
rect 8138 3542 8298 4298
rect 8138 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8298 3542
rect 8138 2758 8298 3514
rect 8138 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8298 2758
rect 8138 1974 8298 2730
rect 8138 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8298 1974
rect 8138 1538 8298 1946
rect 9216 7854 9376 8262
rect 9216 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9376 7854
rect 9216 7070 9376 7826
rect 9216 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9376 7070
rect 9216 6286 9376 7042
rect 9216 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9376 6286
rect 9216 5502 9376 6258
rect 9216 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9376 5502
rect 9216 4718 9376 5474
rect 9216 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9376 4718
rect 9216 3934 9376 4690
rect 9216 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9376 3934
rect 9216 3150 9376 3906
rect 9216 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9376 3150
rect 9216 2366 9376 3122
rect 9216 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9376 2366
rect 9216 1582 9376 2338
rect 9216 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9376 1582
rect 9216 1538 9376 1554
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _083_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7448 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _084_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4984 0 -1 3920
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _085_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4536 0 1 3136
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _086_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2856 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _087_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 -1 3920
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _088_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2800 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _089_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5768 0 1 3920
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _090_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 3136
box -43 -43 1107 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7336 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5712 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _093_
timestamp 1698431365
transform 1 0 7336 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7000 0 -1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _095_
timestamp 1698431365
transform 1 0 7560 0 -1 3136
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_
timestamp 1698431365
transform -1 0 7504 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _097_
timestamp 1698431365
transform -1 0 4592 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4760 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698431365
transform 1 0 4312 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _100_
timestamp 1698431365
transform -1 0 6104 0 1 4704
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5768 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _102_
timestamp 1698431365
transform -1 0 5376 0 1 4704
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1698431365
transform 1 0 4424 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6440 0 -1 6272
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5768 0 1 6272
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _106_
timestamp 1698431365
transform -1 0 5152 0 -1 6272
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698431365
transform 1 0 3752 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _108_
timestamp 1698431365
transform 1 0 4984 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698431365
transform -1 0 7336 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1698431365
transform -1 0 6048 0 1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _111_
timestamp 1698431365
transform -1 0 4592 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698431365
transform 1 0 3976 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _113_
timestamp 1698431365
transform 1 0 4200 0 -1 6272
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _114_
timestamp 1698431365
transform 1 0 5208 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _115_
timestamp 1698431365
transform -1 0 8848 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_
timestamp 1698431365
transform 1 0 6776 0 -1 6272
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _117_
timestamp 1698431365
transform 1 0 6664 0 1 5488
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _118_
timestamp 1698431365
transform 1 0 6440 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _119_
timestamp 1698431365
transform 1 0 7504 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698431365
transform 1 0 3416 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7896 0 -1 5488
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_
timestamp 1698431365
transform -1 0 9072 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _123_
timestamp 1698431365
transform 1 0 4704 0 -1 5488
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6104 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _125_
timestamp 1698431365
transform -1 0 6552 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _126_
timestamp 1698431365
transform 1 0 7056 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _127_
timestamp 1698431365
transform 1 0 6832 0 1 4704
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698431365
transform 1 0 3080 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698431365
transform -1 0 7000 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6552 0 1 3920
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1698431365
transform 1 0 6664 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698431365
transform -1 0 5992 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _134_
timestamp 1698431365
transform -1 0 6832 0 -1 7056
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _135_
timestamp 1698431365
transform 1 0 6664 0 1 6272
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _136_
timestamp 1698431365
transform -1 0 6104 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _137_
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _138_
timestamp 1698431365
transform 1 0 2744 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _139_
timestamp 1698431365
transform 1 0 3248 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2856 0 1 4704
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _141_
timestamp 1698431365
transform 1 0 1344 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _142_
timestamp 1698431365
transform 1 0 2744 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _143_
timestamp 1698431365
transform 1 0 3080 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _144_
timestamp 1698431365
transform -1 0 2744 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _145_
timestamp 1698431365
transform 1 0 1960 0 -1 4704
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _146_
timestamp 1698431365
transform 1 0 1344 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1698431365
transform -1 0 2744 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _148_
timestamp 1698431365
transform -1 0 1960 0 -1 4704
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _149_
timestamp 1698431365
transform -1 0 1568 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698431365
transform -1 0 2408 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _151_
timestamp 1698431365
transform -1 0 1512 0 -1 6272
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1698431365
transform 1 0 1344 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698431365
transform 1 0 2128 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _154_
timestamp 1698431365
transform 1 0 1512 0 -1 6272
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _156_
timestamp 1698431365
transform 1 0 3528 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _157_
timestamp 1698431365
transform 1 0 2968 0 1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698431365
transform -1 0 4984 0 -1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698431365
transform -1 0 3248 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _160_
timestamp 1698431365
transform 1 0 7840 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _161_
timestamp 1698431365
transform 1 0 7168 0 1 6272
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698431365
transform 1 0 6832 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698431365
transform -1 0 7728 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _164_
timestamp 1698431365
transform -1 0 7448 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _166_
timestamp 1698431365
transform 1 0 8624 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4032 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _168_
timestamp 1698431365
transform 1 0 3360 0 1 3920
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7448 0 1 4704
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _170_
timestamp 1698431365
transform 1 0 7392 0 1 3920
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _171_
timestamp 1698431365
transform -1 0 7000 0 -1 3136
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _172_
timestamp 1698431365
transform -1 0 6496 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _173_
timestamp 1698431365
transform 1 0 2744 0 -1 5488
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _174_
timestamp 1698431365
transform 1 0 1008 0 1 3920
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1698431365
transform 1 0 1008 0 1 4704
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1698431365
transform 1 0 1008 0 1 5488
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _177_
timestamp 1698431365
transform 1 0 1008 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1698431365
transform 1 0 2744 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1698431365
transform 1 0 7560 0 1 5488
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1698431365
transform 1 0 6552 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _182_
timestamp 1698431365
transform 1 0 7448 0 1 3136
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6888 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__C
timestamp 1698431365
transform 1 0 3528 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__B
timestamp 1698431365
transform -1 0 7000 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__B
timestamp 1698431365
transform 1 0 8736 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 4480 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1232 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 1232 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 1232 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 1232 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 1120 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 1232 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 8848 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5096 0 -1 5488
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 6048 0 1 5488
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 5712 0 -1 4704
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_28 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_32 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138
timestamp 1698431365
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698431365
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1698431365
transform 1 0 1120 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_12
timestamp 1698431365
transform 1 0 1344 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_44 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_60 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4032 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_68
timestamp 1698431365
transform 1 0 4480 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_150
timestamp 1698431365
transform 1 0 9072 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_43
timestamp 1698431365
transform 1 0 3080 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_75
timestamp 1698431365
transform 1 0 4872 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_91
timestamp 1698431365
transform 1 0 5768 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_99
timestamp 1698431365
transform 1 0 6216 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_103
timestamp 1698431365
transform 1 0 6440 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 6664 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_111
timestamp 1698431365
transform 1 0 6888 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_115
timestamp 1698431365
transform 1 0 7112 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_121
timestamp 1698431365
transform 1 0 7448 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_137
timestamp 1698431365
transform 1 0 8344 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_145
timestamp 1698431365
transform 1 0 8792 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_149
timestamp 1698431365
transform 1 0 9016 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_151
timestamp 1698431365
transform 1 0 9128 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_72
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_80
timestamp 1698431365
transform 1 0 5152 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_146
timestamp 1698431365
transform 1 0 8848 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 9072 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_8
timestamp 1698431365
transform 1 0 1120 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_16
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_66
timestamp 1698431365
transform 1 0 4368 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_68
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_84
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_119
timestamp 1698431365
transform 1 0 7336 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_2
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_10
timestamp 1698431365
transform 1 0 1232 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_16
timestamp 1698431365
transform 1 0 1568 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_24
timestamp 1698431365
transform 1 0 2016 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_28
timestamp 1698431365
transform 1 0 2240 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_59
timestamp 1698431365
transform 1 0 3976 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_61
timestamp 1698431365
transform 1 0 4088 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_150
timestamp 1698431365
transform 1 0 9072 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698431365
transform 1 0 2744 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_45
timestamp 1698431365
transform 1 0 3192 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_47
timestamp 1698431365
transform 1 0 3304 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_119
timestamp 1698431365
transform 1 0 7336 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_149
timestamp 1698431365
transform 1 0 9016 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_151
timestamp 1698431365
transform 1 0 9128 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_8
timestamp 1698431365
transform 1 0 1120 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_12
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_33
timestamp 1698431365
transform 1 0 2520 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_49
timestamp 1698431365
transform 1 0 3416 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_57
timestamp 1698431365
transform 1 0 3864 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_61
timestamp 1698431365
transform 1 0 4088 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_72
timestamp 1698431365
transform 1 0 4704 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_89
timestamp 1698431365
transform 1 0 5656 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_147
timestamp 1698431365
transform 1 0 8904 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_151
timestamp 1698431365
transform 1 0 9128 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_49
timestamp 1698431365
transform 1 0 3416 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_53
timestamp 1698431365
transform 1 0 3640 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_57
timestamp 1698431365
transform 1 0 3864 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 6664 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_109
timestamp 1698431365
transform 1 0 6776 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_8
timestamp 1698431365
transform 1 0 1120 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_16
timestamp 1698431365
transform 1 0 1568 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_24
timestamp 1698431365
transform 1 0 2016 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_66
timestamp 1698431365
transform 1 0 4368 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_150
timestamp 1698431365
transform 1 0 9072 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2
timestamp 1698431365
transform 1 0 784 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_45
timestamp 1698431365
transform 1 0 3192 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_96
timestamp 1698431365
transform 1 0 6048 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_120
timestamp 1698431365
transform 1 0 7392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_122
timestamp 1698431365
transform 1 0 7504 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 784 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_4
timestamp 1698431365
transform 1 0 896 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_25
timestamp 1698431365
transform 1 0 2072 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_32
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_40
timestamp 1698431365
transform 1 0 2912 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_44
timestamp 1698431365
transform 1 0 3136 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_52
timestamp 1698431365
transform 1 0 3584 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_60
timestamp 1698431365
transform 1 0 4032 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_62
timestamp 1698431365
transform 1 0 4144 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_72
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_114
timestamp 1698431365
transform 1 0 7056 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_134
timestamp 1698431365
transform 1 0 8176 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 8400 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2
timestamp 1698431365
transform 1 0 784 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_37
timestamp 1698431365
transform 1 0 2744 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_53
timestamp 1698431365
transform 1 0 3640 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_61
timestamp 1698431365
transform 1 0 4088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_65
timestamp 1698431365
transform 1 0 4312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_73
timestamp 1698431365
transform 1 0 4760 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_75
timestamp 1698431365
transform 1 0 4872 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_97
timestamp 1698431365
transform 1 0 6104 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_114
timestamp 1698431365
transform 1 0 7056 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_8
timestamp 1698431365
transform 1 0 1120 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_16
timestamp 1698431365
transform 1 0 1568 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_24
timestamp 1698431365
transform 1 0 2016 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_28
timestamp 1698431365
transform 1 0 2240 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_30
timestamp 1698431365
transform 1 0 2352 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_61
timestamp 1698431365
transform 1 0 4088 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 4536 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_72
timestamp 1698431365
transform 1 0 4704 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_76
timestamp 1698431365
transform 1 0 4928 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_115
timestamp 1698431365
transform 1 0 7112 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_131
timestamp 1698431365
transform 1 0 8008 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 8456 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 9072 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_2
timestamp 1698431365
transform 1 0 784 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_10
timestamp 1698431365
transform 1 0 1232 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_16
timestamp 1698431365
transform 1 0 1568 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_32
timestamp 1698431365
transform 1 0 2464 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698431365
transform 1 0 2744 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_57
timestamp 1698431365
transform 1 0 3864 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_59
timestamp 1698431365
transform 1 0 3976 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_97
timestamp 1698431365
transform 1 0 6104 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 6664 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_126
timestamp 1698431365
transform 1 0 7728 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_142
timestamp 1698431365
transform 1 0 8624 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_150
timestamp 1698431365
transform 1 0 9072 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 784 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_8
timestamp 1698431365
transform 1 0 1120 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_16
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_32
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_36
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_74
timestamp 1698431365
transform 1 0 4816 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_104
timestamp 1698431365
transform 1 0 6496 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_134
timestamp 1698431365
transform 1 0 8176 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_14
timestamp 1698431365
transform 1 0 1456 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_18
timestamp 1698431365
transform 1 0 1680 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_36
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_70
timestamp 1698431365
transform 1 0 4592 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_104
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_108
timestamp 1698431365
transform 1 0 6720 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_144
timestamp 1698431365
transform 1 0 8736 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 8736 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 784 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 784 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 1120 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform -1 0 9184 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2240 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform 1 0 7728 0 1 6272
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698431365
transform -1 0 8288 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform 1 0 7056 0 -1 3920
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_17 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 9296 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_18
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_19
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 9296 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_20
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 9296 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_21
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 9296 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_22
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 9296 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_23
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 9296 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_24
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 9296 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_25
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 9296 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_26
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 9296 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_27
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 9296 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_28
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 9296 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_29
timestamp 1698431365
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 9296 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_30
timestamp 1698431365
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 9296 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_31
timestamp 1698431365
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 9296 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_32
timestamp 1698431365
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 9296 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_33
timestamp 1698431365
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 9296 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_38
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1698431365
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_40
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_41
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_42
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_43
timestamp 1698431365
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_44
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_45
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_46
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_47
timestamp 1698431365
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_48
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_49
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_50
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_51
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_52
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_53
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_54
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_55
timestamp 1698431365
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_56
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_57
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_58
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_59
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_60
timestamp 1698431365
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_61
timestamp 1698431365
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_62
timestamp 1698431365
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_63
timestamp 1698431365
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_64
timestamp 1698431365
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_65
timestamp 1698431365
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_66
timestamp 1698431365
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_67
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_68
timestamp 1698431365
transform 1 0 2576 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_69
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_70
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_71
timestamp 1698431365
transform 1 0 8288 0 1 7840
box -43 -43 155 435
<< labels >>
flabel metal2 s 2464 9600 2520 10000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 7392 9600 7448 10000 0 FreeSans 224 90 0 0 reset
port 1 nsew signal input
flabel metal3 s 0 3024 400 3080 0 FreeSans 224 0 0 0 rle1__input_r[0]
port 2 nsew signal input
flabel metal3 s 0 4256 400 4312 0 FreeSans 224 0 0 0 rle1__input_r[1]
port 3 nsew signal input
flabel metal3 s 0 5488 400 5544 0 FreeSans 224 0 0 0 rle1__input_r[2]
port 4 nsew signal input
flabel metal3 s 0 6720 400 6776 0 FreeSans 224 0 0 0 rle1__input_r[3]
port 5 nsew signal input
flabel metal3 s 0 7952 400 8008 0 FreeSans 224 0 0 0 rle1__input_r[4]
port 6 nsew signal input
flabel metal3 s 0 9184 400 9240 0 FreeSans 224 0 0 0 rle1__input_r[5]
port 7 nsew signal input
flabel metal3 s 0 560 400 616 0 FreeSans 224 0 0 0 rle1__input_r_rdy
port 8 nsew signal tristate
flabel metal3 s 0 1792 400 1848 0 FreeSans 224 0 0 0 rle1__input_r_vld
port 9 nsew signal input
flabel metal3 s 9600 6160 10000 6216 0 FreeSans 224 0 0 0 rle1__output_s[0]
port 10 nsew signal tristate
flabel metal3 s 9600 8624 10000 8680 0 FreeSans 224 0 0 0 rle1__output_s[1]
port 11 nsew signal tristate
flabel metal3 s 9600 1232 10000 1288 0 FreeSans 224 0 0 0 rle1__output_s_rdy
port 12 nsew signal input
flabel metal3 s 9600 3696 10000 3752 0 FreeSans 224 0 0 0 rle1__output_s_vld
port 13 nsew signal tristate
flabel metal4 s 1670 1538 1830 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 3826 1538 3986 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 5982 1538 6142 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 8138 1538 8298 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 2748 1538 2908 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 4904 1538 5064 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 7060 1538 7220 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 9216 1538 9376 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
rlabel metal1 4984 8232 4984 8232 0 vdd
rlabel via1 5024 7840 5024 7840 0 vss
rlabel metal2 5124 7084 5124 7084 0 _000_
rlabel metal2 3836 4200 3836 4200 0 _001_
rlabel metal2 7952 4956 7952 4956 0 _002_
rlabel metal3 7644 4172 7644 4172 0 _003_
rlabel metal2 6524 3192 6524 3192 0 _004_
rlabel metal2 5908 7364 5908 7364 0 _005_
rlabel metal2 3108 5012 3108 5012 0 _006_
rlabel metal3 1792 4396 1792 4396 0 _007_
rlabel metal2 1484 4732 1484 4732 0 _008_
rlabel metal2 1372 5880 1372 5880 0 _009_
rlabel metal2 1484 6300 1484 6300 0 _010_
rlabel metal2 3220 7364 3220 7364 0 _011_
rlabel metal2 3220 3416 3220 3416 0 _012_
rlabel metal3 7756 5628 7756 5628 0 _013_
rlabel metal2 7308 7448 7308 7448 0 _014_
rlabel metal2 7924 3500 7924 3500 0 _015_
rlabel metal2 1512 3836 1512 3836 0 _016_
rlabel metal2 2324 5656 2324 5656 0 _017_
rlabel metal2 3220 4424 3220 4424 0 _018_
rlabel metal2 1988 6132 1988 6132 0 _019_
rlabel metal2 1708 4732 1708 4732 0 _020_
rlabel metal2 1652 4704 1652 4704 0 _021_
rlabel metal2 1316 6440 1316 6440 0 _022_
rlabel metal2 2156 5404 2156 5404 0 _023_
rlabel metal2 1708 6356 1708 6356 0 _024_
rlabel metal2 2212 6076 2212 6076 0 _025_
rlabel metal2 3164 7448 3164 7448 0 _026_
rlabel metal3 3472 7252 3472 7252 0 _027_
rlabel metal2 3220 3752 3220 3752 0 _028_
rlabel metal2 7980 6328 7980 6328 0 _029_
rlabel metal2 7168 6972 7168 6972 0 _030_
rlabel metal2 7420 7196 7420 7196 0 _031_
rlabel metal2 8876 4144 8876 4144 0 _032_
rlabel metal2 6188 2996 6188 2996 0 _033_
rlabel metal3 4816 3836 4816 3836 0 _034_
rlabel metal2 4956 3584 4956 3584 0 _035_
rlabel metal2 2996 3192 2996 3192 0 _036_
rlabel metal3 3052 3836 3052 3836 0 _037_
rlabel metal2 5796 3108 5796 3108 0 _038_
rlabel metal2 7196 3388 7196 3388 0 _039_
rlabel metal2 7644 7056 7644 7056 0 _040_
rlabel metal2 5376 6972 5376 6972 0 _041_
rlabel metal2 8204 3136 8204 3136 0 _042_
rlabel metal3 8204 2940 8204 2940 0 _043_
rlabel metal2 7756 3626 7756 3626 0 _044_
rlabel metal3 4676 6188 4676 6188 0 _045_
rlabel metal3 5152 4900 5152 4900 0 _046_
rlabel metal2 4872 4620 4872 4620 0 _047_
rlabel metal2 6188 4704 6188 4704 0 _048_
rlabel metal2 5628 5516 5628 5516 0 _049_
rlabel metal2 6860 5992 6860 5992 0 _050_
rlabel via2 4900 6132 4900 6132 0 _051_
rlabel metal2 6356 6244 6356 6244 0 _052_
rlabel metal3 5516 6076 5516 6076 0 _053_
rlabel metal2 5656 6412 5656 6412 0 _054_
rlabel metal2 4788 6524 4788 6524 0 _055_
rlabel metal2 2940 3864 2940 3864 0 _056_
rlabel metal3 6916 3836 6916 3836 0 _057_
rlabel metal2 5656 4396 5656 4396 0 _058_
rlabel metal2 4396 4956 4396 4956 0 _059_
rlabel metal2 4312 6076 4312 6076 0 _060_
rlabel metal2 5236 5040 5236 5040 0 _061_
rlabel metal2 8568 5292 8568 5292 0 _062_
rlabel metal2 6944 5628 6944 5628 0 _063_
rlabel metal3 7560 5292 7560 5292 0 _064_
rlabel metal3 7140 5964 7140 5964 0 _065_
rlabel metal2 7924 5432 7924 5432 0 _066_
rlabel metal2 3668 6692 3668 6692 0 _067_
rlabel metal2 7364 5040 7364 5040 0 _068_
rlabel metal2 6328 4116 6328 4116 0 _069_
rlabel metal2 7028 4956 7028 4956 0 _070_
rlabel metal2 6412 5292 6412 5292 0 _071_
rlabel metal2 6916 5208 6916 5208 0 _072_
rlabel metal2 3332 7084 3332 7084 0 _073_
rlabel metal2 6804 4144 6804 4144 0 _074_
rlabel metal3 6748 3332 6748 3332 0 _075_
rlabel metal2 5768 6972 5768 6972 0 _076_
rlabel metal2 6832 6356 6832 6356 0 _077_
rlabel metal2 6804 6860 6804 6860 0 _078_
rlabel metal3 6496 6580 6496 6580 0 _079_
rlabel metal3 2268 3332 2268 3332 0 _080_
rlabel metal2 1512 6076 1512 6076 0 _081_
rlabel metal2 3220 5068 3220 5068 0 _082_
rlabel metal2 2492 8589 2492 8589 0 clk
rlabel metal2 5852 5516 5852 5516 0 clknet_0_clk
rlabel metal3 3164 3612 3164 3612 0 clknet_1_0__leaf_clk
rlabel metal2 7532 3136 7532 3136 0 clknet_1_1__leaf_clk
rlabel metal2 3892 6916 3892 6916 0 net1
rlabel metal2 2436 2716 2436 2716 0 net10
rlabel metal2 8036 5936 8036 5936 0 net11
rlabel metal2 8092 7812 8092 7812 0 net12
rlabel metal2 8988 3416 8988 3416 0 net13
rlabel metal2 1036 3304 1036 3304 0 net2
rlabel metal2 1428 3892 1428 3892 0 net3
rlabel metal3 1232 5236 1232 5236 0 net4
rlabel metal2 1260 6916 1260 6916 0 net5
rlabel metal2 1428 7420 1428 7420 0 net6
rlabel metal2 1428 7812 1428 7812 0 net7
rlabel metal2 1036 2408 1036 2408 0 net8
rlabel metal2 7420 2856 7420 2856 0 net9
rlabel metal3 8008 8036 8008 8036 0 reset
rlabel metal2 868 3164 868 3164 0 rle1__input_r[0]
rlabel metal2 868 4396 868 4396 0 rle1__input_r[1]
rlabel metal2 868 5432 868 5432 0 rle1__input_r[2]
rlabel metal2 868 6804 868 6804 0 rle1__input_r[3]
rlabel metal3 623 7980 623 7980 0 rle1__input_r[4]
rlabel metal2 1204 8624 1204 8624 0 rle1__input_r[5]
rlabel metal3 427 588 427 588 0 rle1__input_r_rdy
rlabel metal2 868 1988 868 1988 0 rle1__input_r_vld
rlabel metal2 8988 6356 8988 6356 0 rle1__output_s[0]
rlabel metal3 8561 8652 8561 8652 0 rle1__output_s[1]
rlabel metal2 9100 1484 9100 1484 0 rle1__output_s_rdy
rlabel metal2 8316 3696 8316 3696 0 rle1__output_s_vld
rlabel metal2 5852 7028 5852 7028 0 rle1_dec_0.____state_0
rlabel metal3 4592 4172 4592 4172 0 rle1_dec_0.____state_1\[0\]
rlabel metal2 5124 3724 5124 3724 0 rle1_dec_0.____state_1\[1\]
rlabel metal3 7000 3724 7000 3724 0 rle1_dec_0.____state_1\[2\]
rlabel metal2 5656 4060 5656 4060 0 rle1_dec_0.____state_1\[3\]
rlabel metal2 5572 6748 5572 6748 0 rle1_dec_0.____state_2
rlabel metal2 3500 6132 3500 6132 0 rle1_dec_0.__rle1__input_r_reg\[0\]
rlabel metal3 2940 4508 2940 4508 0 rle1_dec_0.__rle1__input_r_reg\[1\]
rlabel metal2 2548 4928 2548 4928 0 rle1_dec_0.__rle1__input_r_reg\[2\]
rlabel metal2 2212 5264 2212 5264 0 rle1_dec_0.__rle1__input_r_reg\[3\]
rlabel metal2 2380 5992 2380 5992 0 rle1_dec_0.__rle1__input_r_reg\[4\]
rlabel metal2 3780 7280 3780 7280 0 rle1_dec_0.__rle1__input_r_reg\[5\]
rlabel metal2 3780 3696 3780 3696 0 rle1_dec_0.__rle1__input_r_valid_reg
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
