magic
tech gf180mcuD
magscale 1 5
timestamp 1702516937
<< metal1 >>
rect 672 8245 9296 8262
rect 672 8219 1685 8245
rect 1711 8219 1737 8245
rect 1763 8219 1789 8245
rect 1815 8219 3841 8245
rect 3867 8219 3893 8245
rect 3919 8219 3945 8245
rect 3971 8219 5997 8245
rect 6023 8219 6049 8245
rect 6075 8219 6101 8245
rect 6127 8219 8153 8245
rect 8179 8219 8205 8245
rect 8231 8219 8257 8245
rect 8283 8219 9296 8245
rect 672 8202 9296 8219
rect 1247 8105 1273 8111
rect 1247 8073 1273 8079
rect 8863 8105 8889 8111
rect 8863 8073 8889 8079
rect 855 8049 881 8055
rect 8185 8023 8191 8049
rect 8217 8023 8223 8049
rect 8577 8023 8583 8049
rect 8609 8023 8615 8049
rect 855 8017 881 8023
rect 6119 7993 6145 7999
rect 7401 7967 7407 7993
rect 7433 7967 7439 7993
rect 6119 7961 6145 7967
rect 1023 7937 1049 7943
rect 1023 7905 1049 7911
rect 6287 7937 6313 7943
rect 6287 7905 6313 7911
rect 8471 7937 8497 7943
rect 8471 7905 8497 7911
rect 672 7853 9376 7870
rect 672 7827 2763 7853
rect 2789 7827 2815 7853
rect 2841 7827 2867 7853
rect 2893 7827 4919 7853
rect 4945 7827 4971 7853
rect 4997 7827 5023 7853
rect 5049 7827 7075 7853
rect 7101 7827 7127 7853
rect 7153 7827 7179 7853
rect 7205 7827 9231 7853
rect 9257 7827 9283 7853
rect 9309 7827 9335 7853
rect 9361 7827 9376 7853
rect 672 7810 9376 7827
rect 7911 7769 7937 7775
rect 7911 7737 7937 7743
rect 8807 7769 8833 7775
rect 8807 7737 8833 7743
rect 3033 7631 3039 7657
rect 3065 7631 3071 7657
rect 3425 7631 3431 7657
rect 3457 7631 3463 7657
rect 6897 7631 6903 7657
rect 6929 7631 6935 7657
rect 8409 7631 8415 7657
rect 8441 7631 8447 7657
rect 4887 7601 4913 7607
rect 4489 7575 4495 7601
rect 4521 7575 4527 7601
rect 5441 7575 5447 7601
rect 5473 7575 5479 7601
rect 6505 7575 6511 7601
rect 6537 7575 6543 7601
rect 8801 7575 8807 7601
rect 8833 7575 8839 7601
rect 4887 7569 4913 7575
rect 8695 7545 8721 7551
rect 8695 7513 8721 7519
rect 672 7461 9296 7478
rect 672 7435 1685 7461
rect 1711 7435 1737 7461
rect 1763 7435 1789 7461
rect 1815 7435 3841 7461
rect 3867 7435 3893 7461
rect 3919 7435 3945 7461
rect 3971 7435 5997 7461
rect 6023 7435 6049 7461
rect 6075 7435 6101 7461
rect 6127 7435 8153 7461
rect 8179 7435 8205 7461
rect 8231 7435 8257 7461
rect 8283 7435 9296 7461
rect 672 7418 9296 7435
rect 5951 7377 5977 7383
rect 5951 7345 5977 7351
rect 4327 7321 4353 7327
rect 4327 7289 4353 7295
rect 6399 7321 6425 7327
rect 9025 7295 9031 7321
rect 9057 7295 9063 7321
rect 6399 7289 6425 7295
rect 4551 7265 4577 7271
rect 4551 7233 4577 7239
rect 4943 7265 4969 7271
rect 4943 7233 4969 7239
rect 5111 7265 5137 7271
rect 5895 7265 5921 7271
rect 5329 7239 5335 7265
rect 5361 7239 5367 7265
rect 5111 7233 5137 7239
rect 5895 7233 5921 7239
rect 7239 7265 7265 7271
rect 7289 7239 7295 7265
rect 7321 7239 7327 7265
rect 7569 7239 7575 7265
rect 7601 7239 7607 7265
rect 7239 7233 7265 7239
rect 4775 7209 4801 7215
rect 5559 7209 5585 7215
rect 4881 7183 4887 7209
rect 4913 7183 4919 7209
rect 4775 7177 4801 7183
rect 5559 7177 5585 7183
rect 6231 7209 6257 7215
rect 6231 7177 6257 7183
rect 6455 7209 6481 7215
rect 6455 7177 6481 7183
rect 7015 7209 7041 7215
rect 7121 7183 7127 7209
rect 7153 7183 7159 7209
rect 7961 7183 7967 7209
rect 7993 7183 7999 7209
rect 7015 7177 7041 7183
rect 3935 7153 3961 7159
rect 4439 7153 4465 7159
rect 4097 7127 4103 7153
rect 4129 7127 4135 7153
rect 3935 7121 3961 7127
rect 4439 7121 4465 7127
rect 5167 7153 5193 7159
rect 5167 7121 5193 7127
rect 5615 7153 5641 7159
rect 5615 7121 5641 7127
rect 5671 7153 5697 7159
rect 5671 7121 5697 7127
rect 5727 7153 5753 7159
rect 5727 7121 5753 7127
rect 6007 7153 6033 7159
rect 6007 7121 6033 7127
rect 6119 7153 6145 7159
rect 6119 7121 6145 7127
rect 7407 7153 7433 7159
rect 7407 7121 7433 7127
rect 672 7069 9376 7086
rect 672 7043 2763 7069
rect 2789 7043 2815 7069
rect 2841 7043 2867 7069
rect 2893 7043 4919 7069
rect 4945 7043 4971 7069
rect 4997 7043 5023 7069
rect 5049 7043 7075 7069
rect 7101 7043 7127 7069
rect 7153 7043 7179 7069
rect 7205 7043 9231 7069
rect 9257 7043 9283 7069
rect 9309 7043 9335 7069
rect 9361 7043 9376 7069
rect 672 7026 9376 7043
rect 4551 6985 4577 6991
rect 4551 6953 4577 6959
rect 6063 6985 6089 6991
rect 6063 6953 6089 6959
rect 6679 6985 6705 6991
rect 6679 6953 6705 6959
rect 6903 6985 6929 6991
rect 6903 6953 6929 6959
rect 8751 6985 8777 6991
rect 8751 6953 8777 6959
rect 4495 6929 4521 6935
rect 4495 6897 4521 6903
rect 4775 6929 4801 6935
rect 4775 6897 4801 6903
rect 4887 6873 4913 6879
rect 2641 6847 2647 6873
rect 2673 6847 2679 6873
rect 4265 6847 4271 6873
rect 4297 6847 4303 6873
rect 4377 6847 4383 6873
rect 4409 6847 4415 6873
rect 4887 6841 4913 6847
rect 4999 6873 5025 6879
rect 6175 6873 6201 6879
rect 5833 6847 5839 6873
rect 5865 6847 5871 6873
rect 5945 6847 5951 6873
rect 5977 6847 5983 6873
rect 4999 6841 5025 6847
rect 6175 6841 6201 6847
rect 6287 6873 6313 6879
rect 6287 6841 6313 6847
rect 6399 6873 6425 6879
rect 6959 6873 6985 6879
rect 6561 6847 6567 6873
rect 6593 6847 6599 6873
rect 8409 6847 8415 6873
rect 8441 6847 8447 6873
rect 8857 6847 8863 6873
rect 8889 6847 8895 6873
rect 6399 6841 6425 6847
rect 6959 6841 6985 6847
rect 6511 6817 6537 6823
rect 2977 6791 2983 6817
rect 3009 6791 3015 6817
rect 4041 6791 4047 6817
rect 4073 6791 4079 6817
rect 6511 6785 6537 6791
rect 5111 6761 5137 6767
rect 5111 6729 5137 6735
rect 5335 6761 5361 6767
rect 5335 6729 5361 6735
rect 6063 6761 6089 6767
rect 6063 6729 6089 6735
rect 6903 6761 6929 6767
rect 6903 6729 6929 6735
rect 7911 6761 7937 6767
rect 7911 6729 7937 6735
rect 8695 6761 8721 6767
rect 8695 6729 8721 6735
rect 672 6677 9296 6694
rect 672 6651 1685 6677
rect 1711 6651 1737 6677
rect 1763 6651 1789 6677
rect 1815 6651 3841 6677
rect 3867 6651 3893 6677
rect 3919 6651 3945 6677
rect 3971 6651 5997 6677
rect 6023 6651 6049 6677
rect 6075 6651 6101 6677
rect 6127 6651 8153 6677
rect 8179 6651 8205 6677
rect 8231 6651 8257 6677
rect 8283 6651 9296 6677
rect 672 6634 9296 6651
rect 5055 6593 5081 6599
rect 5055 6561 5081 6567
rect 5167 6593 5193 6599
rect 5167 6561 5193 6567
rect 5783 6593 5809 6599
rect 5783 6561 5809 6567
rect 5335 6537 5361 6543
rect 4041 6511 4047 6537
rect 4073 6511 4079 6537
rect 8017 6511 8023 6537
rect 8049 6511 8055 6537
rect 9081 6511 9087 6537
rect 9113 6511 9119 6537
rect 5335 6505 5361 6511
rect 5279 6481 5305 6487
rect 4209 6455 4215 6481
rect 4241 6455 4247 6481
rect 4713 6455 4719 6481
rect 4745 6455 4751 6481
rect 5279 6449 5305 6455
rect 5671 6481 5697 6487
rect 5889 6455 5895 6481
rect 5921 6455 5927 6481
rect 6001 6455 6007 6481
rect 6033 6455 6039 6481
rect 7009 6455 7015 6481
rect 7041 6455 7047 6481
rect 7625 6455 7631 6481
rect 7657 6455 7663 6481
rect 5671 6449 5697 6455
rect 855 6425 881 6431
rect 855 6393 881 6399
rect 4439 6425 4465 6431
rect 4439 6393 4465 6399
rect 4607 6425 4633 6431
rect 4607 6393 4633 6399
rect 5559 6425 5585 6431
rect 5559 6393 5585 6399
rect 6175 6425 6201 6431
rect 6175 6393 6201 6399
rect 6343 6425 6369 6431
rect 6343 6393 6369 6399
rect 7295 6425 7321 6431
rect 7295 6393 7321 6399
rect 1023 6369 1049 6375
rect 1023 6337 1049 6343
rect 1247 6369 1273 6375
rect 1247 6337 1273 6343
rect 5335 6369 5361 6375
rect 5335 6337 5361 6343
rect 5783 6369 5809 6375
rect 5783 6337 5809 6343
rect 7127 6369 7153 6375
rect 7127 6337 7153 6343
rect 7463 6369 7489 6375
rect 7463 6337 7489 6343
rect 672 6285 9376 6302
rect 672 6259 2763 6285
rect 2789 6259 2815 6285
rect 2841 6259 2867 6285
rect 2893 6259 4919 6285
rect 4945 6259 4971 6285
rect 4997 6259 5023 6285
rect 5049 6259 7075 6285
rect 7101 6259 7127 6285
rect 7153 6259 7179 6285
rect 7205 6259 9231 6285
rect 9257 6259 9283 6285
rect 9309 6259 9335 6285
rect 9361 6259 9376 6285
rect 672 6242 9376 6259
rect 3599 6201 3625 6207
rect 3599 6169 3625 6175
rect 3823 6201 3849 6207
rect 3823 6169 3849 6175
rect 4047 6201 4073 6207
rect 4047 6169 4073 6175
rect 4831 6201 4857 6207
rect 5217 6175 5223 6201
rect 5249 6175 5255 6201
rect 4831 6169 4857 6175
rect 4271 6145 4297 6151
rect 4271 6113 4297 6119
rect 4495 6145 4521 6151
rect 5951 6145 5977 6151
rect 5721 6119 5727 6145
rect 5753 6119 5759 6145
rect 4495 6113 4521 6119
rect 5951 6113 5977 6119
rect 6791 6145 6817 6151
rect 6791 6113 6817 6119
rect 6959 6145 6985 6151
rect 6959 6113 6985 6119
rect 3991 6089 4017 6095
rect 4999 6089 5025 6095
rect 1969 6063 1975 6089
rect 2001 6063 2007 6089
rect 4377 6063 4383 6089
rect 4409 6063 4415 6089
rect 3991 6057 4017 6063
rect 4999 6057 5025 6063
rect 5167 6089 5193 6095
rect 5559 6089 5585 6095
rect 8639 6089 8665 6095
rect 5329 6063 5335 6089
rect 5361 6063 5367 6089
rect 6393 6063 6399 6089
rect 6425 6063 6431 6089
rect 8353 6063 8359 6089
rect 8385 6063 8391 6089
rect 5167 6057 5193 6063
rect 5559 6057 5585 6063
rect 8639 6057 8665 6063
rect 8863 6089 8889 6095
rect 8863 6057 8889 6063
rect 8919 6089 8945 6095
rect 8919 6057 8945 6063
rect 6287 6033 6313 6039
rect 2305 6007 2311 6033
rect 2337 6007 2343 6033
rect 3369 6007 3375 6033
rect 3401 6007 3407 6033
rect 6287 6001 6313 6007
rect 8751 6033 8777 6039
rect 8751 6001 8777 6007
rect 4047 5977 4073 5983
rect 4047 5945 4073 5951
rect 4551 5977 4577 5983
rect 5895 5977 5921 5983
rect 5273 5951 5279 5977
rect 5305 5951 5311 5977
rect 4551 5945 4577 5951
rect 5895 5945 5921 5951
rect 6063 5977 6089 5983
rect 6063 5945 6089 5951
rect 6231 5977 6257 5983
rect 6231 5945 6257 5951
rect 7911 5977 7937 5983
rect 7911 5945 7937 5951
rect 672 5893 9296 5910
rect 672 5867 1685 5893
rect 1711 5867 1737 5893
rect 1763 5867 1789 5893
rect 1815 5867 3841 5893
rect 3867 5867 3893 5893
rect 3919 5867 3945 5893
rect 3971 5867 5997 5893
rect 6023 5867 6049 5893
rect 6075 5867 6101 5893
rect 6127 5867 8153 5893
rect 8179 5867 8205 5893
rect 8231 5867 8257 5893
rect 8283 5867 9296 5893
rect 672 5850 9296 5867
rect 5727 5809 5753 5815
rect 5161 5783 5167 5809
rect 5193 5783 5199 5809
rect 5727 5777 5753 5783
rect 1415 5753 1441 5759
rect 1415 5721 1441 5727
rect 1695 5753 1721 5759
rect 4943 5753 4969 5759
rect 4265 5727 4271 5753
rect 4297 5727 4303 5753
rect 1695 5721 1721 5727
rect 4943 5721 4969 5727
rect 7295 5753 7321 5759
rect 8017 5727 8023 5753
rect 8049 5727 8055 5753
rect 9081 5727 9087 5753
rect 9113 5727 9119 5753
rect 7295 5721 7321 5727
rect 1471 5697 1497 5703
rect 4607 5697 4633 5703
rect 2809 5671 2815 5697
rect 2841 5671 2847 5697
rect 1471 5665 1497 5671
rect 4607 5665 4633 5671
rect 4887 5697 4913 5703
rect 6063 5697 6089 5703
rect 4993 5671 4999 5697
rect 5025 5671 5031 5697
rect 5161 5671 5167 5697
rect 5193 5671 5199 5697
rect 6337 5671 6343 5697
rect 6369 5671 6375 5697
rect 6841 5671 6847 5697
rect 6873 5671 6879 5697
rect 7177 5671 7183 5697
rect 7209 5671 7215 5697
rect 7345 5671 7351 5697
rect 7377 5671 7383 5697
rect 7625 5671 7631 5697
rect 7657 5671 7663 5697
rect 4887 5665 4913 5671
rect 6063 5665 6089 5671
rect 5895 5641 5921 5647
rect 7071 5641 7097 5647
rect 3201 5615 3207 5641
rect 3233 5615 3239 5641
rect 6729 5615 6735 5641
rect 6761 5615 6767 5641
rect 5895 5609 5921 5615
rect 7071 5609 7097 5615
rect 1639 5585 1665 5591
rect 5615 5585 5641 5591
rect 4433 5559 4439 5585
rect 4465 5559 4471 5585
rect 1639 5553 1665 5559
rect 5615 5553 5641 5559
rect 5671 5585 5697 5591
rect 7463 5585 7489 5591
rect 6225 5559 6231 5585
rect 6257 5559 6263 5585
rect 5671 5553 5697 5559
rect 7463 5553 7489 5559
rect 672 5501 9376 5518
rect 672 5475 2763 5501
rect 2789 5475 2815 5501
rect 2841 5475 2867 5501
rect 2893 5475 4919 5501
rect 4945 5475 4971 5501
rect 4997 5475 5023 5501
rect 5049 5475 7075 5501
rect 7101 5475 7127 5501
rect 7153 5475 7179 5501
rect 7205 5475 9231 5501
rect 9257 5475 9283 5501
rect 9309 5475 9335 5501
rect 9361 5475 9376 5501
rect 672 5458 9376 5475
rect 2535 5417 2561 5423
rect 1465 5391 1471 5417
rect 1497 5391 1503 5417
rect 2535 5385 2561 5391
rect 2815 5417 2841 5423
rect 2815 5385 2841 5391
rect 3151 5417 3177 5423
rect 3151 5385 3177 5391
rect 7911 5417 7937 5423
rect 7911 5385 7937 5391
rect 8751 5417 8777 5423
rect 8751 5385 8777 5391
rect 8863 5417 8889 5423
rect 8863 5385 8889 5391
rect 2759 5361 2785 5367
rect 4775 5361 4801 5367
rect 1409 5335 1415 5361
rect 1441 5335 1447 5361
rect 4265 5335 4271 5361
rect 4297 5335 4303 5361
rect 2759 5329 2785 5335
rect 4775 5329 4801 5335
rect 4831 5361 4857 5367
rect 4831 5329 4857 5335
rect 7855 5361 7881 5367
rect 7855 5329 7881 5335
rect 8191 5361 8217 5367
rect 8191 5329 8217 5335
rect 1303 5305 1329 5311
rect 2983 5305 3009 5311
rect 1633 5279 1639 5305
rect 1665 5279 1671 5305
rect 1303 5273 1329 5279
rect 2983 5273 3009 5279
rect 3207 5305 3233 5311
rect 3207 5273 3233 5279
rect 3319 5305 3345 5311
rect 3319 5273 3345 5279
rect 3487 5305 3513 5311
rect 3487 5273 3513 5279
rect 3599 5305 3625 5311
rect 3599 5273 3625 5279
rect 3767 5305 3793 5311
rect 4943 5305 4969 5311
rect 8135 5305 8161 5311
rect 3929 5279 3935 5305
rect 3961 5279 3967 5305
rect 4489 5279 4495 5305
rect 4521 5279 4527 5305
rect 5105 5279 5111 5305
rect 5137 5279 5143 5305
rect 3767 5273 3793 5279
rect 4943 5273 4969 5279
rect 8135 5273 8161 5279
rect 8303 5305 8329 5311
rect 8303 5273 8329 5279
rect 8695 5305 8721 5311
rect 8695 5273 8721 5279
rect 2871 5249 2897 5255
rect 2871 5217 2897 5223
rect 3711 5249 3737 5255
rect 9031 5249 9057 5255
rect 4433 5223 4439 5249
rect 4465 5223 4471 5249
rect 6169 5223 6175 5249
rect 6201 5223 6207 5249
rect 3711 5217 3737 5223
rect 9031 5217 9057 5223
rect 7911 5193 7937 5199
rect 1577 5167 1583 5193
rect 1609 5167 1615 5193
rect 7911 5161 7937 5167
rect 672 5109 9296 5126
rect 672 5083 1685 5109
rect 1711 5083 1737 5109
rect 1763 5083 1789 5109
rect 1815 5083 3841 5109
rect 3867 5083 3893 5109
rect 3919 5083 3945 5109
rect 3971 5083 5997 5109
rect 6023 5083 6049 5109
rect 6075 5083 6101 5109
rect 6127 5083 8153 5109
rect 8179 5083 8205 5109
rect 8231 5083 8257 5109
rect 8283 5083 9296 5109
rect 672 5066 9296 5083
rect 6225 4999 6231 5025
rect 6257 4999 6263 5025
rect 1465 4943 1471 4969
rect 1497 4943 1503 4969
rect 2529 4943 2535 4969
rect 2561 4943 2567 4969
rect 3649 4943 3655 4969
rect 3681 4943 3687 4969
rect 8969 4943 8975 4969
rect 9001 4943 9007 4969
rect 5951 4913 5977 4919
rect 7127 4913 7153 4919
rect 1129 4887 1135 4913
rect 1161 4887 1167 4913
rect 5721 4887 5727 4913
rect 5753 4887 5759 4913
rect 6337 4887 6343 4913
rect 6369 4887 6375 4913
rect 6841 4887 6847 4913
rect 6873 4887 6879 4913
rect 7569 4887 7575 4913
rect 7601 4887 7607 4913
rect 5951 4881 5977 4887
rect 7127 4881 7153 4887
rect 6057 4831 6063 4857
rect 6089 4831 6095 4857
rect 7289 4831 7295 4857
rect 7321 4831 7327 4857
rect 7905 4831 7911 4857
rect 7937 4831 7943 4857
rect 2983 4801 3009 4807
rect 2983 4769 3009 4775
rect 6343 4801 6369 4807
rect 6953 4775 6959 4801
rect 6985 4775 6991 4801
rect 6343 4769 6369 4775
rect 672 4717 9376 4734
rect 672 4691 2763 4717
rect 2789 4691 2815 4717
rect 2841 4691 2867 4717
rect 2893 4691 4919 4717
rect 4945 4691 4971 4717
rect 4997 4691 5023 4717
rect 5049 4691 7075 4717
rect 7101 4691 7127 4717
rect 7153 4691 7179 4717
rect 7205 4691 9231 4717
rect 9257 4691 9283 4717
rect 9309 4691 9335 4717
rect 9361 4691 9376 4717
rect 672 4674 9376 4691
rect 2647 4633 2673 4639
rect 2647 4601 2673 4607
rect 4831 4633 4857 4639
rect 4831 4601 4857 4607
rect 8751 4633 8777 4639
rect 8751 4601 8777 4607
rect 2759 4577 2785 4583
rect 4775 4577 4801 4583
rect 3369 4551 3375 4577
rect 3401 4551 3407 4577
rect 2759 4545 2785 4551
rect 4775 4545 4801 4551
rect 5615 4577 5641 4583
rect 8695 4577 8721 4583
rect 7569 4551 7575 4577
rect 7601 4551 7607 4577
rect 5615 4545 5641 4551
rect 8695 4545 8721 4551
rect 8975 4577 9001 4583
rect 8975 4545 9001 4551
rect 2815 4521 2841 4527
rect 8863 4521 8889 4527
rect 1129 4495 1135 4521
rect 1161 4495 1167 4521
rect 3033 4495 3039 4521
rect 3065 4495 3071 4521
rect 5329 4495 5335 4521
rect 5361 4495 5367 4521
rect 5777 4495 5783 4521
rect 5809 4495 5815 4521
rect 2815 4489 2841 4495
rect 8863 4489 8889 4495
rect 911 4465 937 4471
rect 1465 4439 1471 4465
rect 1497 4439 1503 4465
rect 2529 4439 2535 4465
rect 2561 4439 2567 4465
rect 4433 4439 4439 4465
rect 4465 4439 4471 4465
rect 5385 4439 5391 4465
rect 5417 4439 5423 4465
rect 911 4433 937 4439
rect 4831 4409 4857 4415
rect 4831 4377 4857 4383
rect 672 4325 9296 4342
rect 672 4299 1685 4325
rect 1711 4299 1737 4325
rect 1763 4299 1789 4325
rect 1815 4299 3841 4325
rect 3867 4299 3893 4325
rect 3919 4299 3945 4325
rect 3971 4299 5997 4325
rect 6023 4299 6049 4325
rect 6075 4299 6101 4325
rect 6127 4299 8153 4325
rect 8179 4299 8205 4325
rect 8231 4299 8257 4325
rect 8283 4299 9296 4325
rect 672 4282 9296 4299
rect 5951 4241 5977 4247
rect 1577 4215 1583 4241
rect 1609 4215 1615 4241
rect 5951 4209 5977 4215
rect 1919 4185 1945 4191
rect 1919 4153 1945 4159
rect 2871 4185 2897 4191
rect 2871 4153 2897 4159
rect 3711 4185 3737 4191
rect 3711 4153 3737 4159
rect 4551 4185 4577 4191
rect 4551 4153 4577 4159
rect 6735 4185 6761 4191
rect 9081 4159 9087 4185
rect 9113 4159 9119 4185
rect 6735 4153 6761 4159
rect 1975 4129 2001 4135
rect 905 4103 911 4129
rect 937 4103 943 4129
rect 1409 4103 1415 4129
rect 1441 4103 1447 4129
rect 1577 4103 1583 4129
rect 1609 4103 1615 4129
rect 1975 4097 2001 4103
rect 2143 4129 2169 4135
rect 6847 4129 6873 4135
rect 5217 4103 5223 4129
rect 5249 4103 5255 4129
rect 5385 4103 5391 4129
rect 5417 4103 5423 4129
rect 7233 4103 7239 4129
rect 7265 4103 7271 4129
rect 7681 4103 7687 4129
rect 7713 4103 7719 4129
rect 2143 4097 2169 4103
rect 6847 4097 6873 4103
rect 1303 4073 1329 4079
rect 1303 4041 1329 4047
rect 1863 4073 1889 4079
rect 5895 4073 5921 4079
rect 4937 4047 4943 4073
rect 4969 4047 4975 4073
rect 1863 4041 1889 4047
rect 5895 4041 5921 4047
rect 6287 4073 6313 4079
rect 6287 4041 6313 4047
rect 6399 4073 6425 4079
rect 8017 4047 8023 4073
rect 8049 4047 8055 4073
rect 6399 4041 6425 4047
rect 1023 4017 1049 4023
rect 3655 4017 3681 4023
rect 1465 3991 1471 4017
rect 1497 3991 1503 4017
rect 1023 3985 1049 3991
rect 3655 3985 3681 3991
rect 3767 4017 3793 4023
rect 3767 3985 3793 3991
rect 3879 4017 3905 4023
rect 3879 3985 3905 3991
rect 6343 4017 6369 4023
rect 7009 3991 7015 4017
rect 7041 3991 7047 4017
rect 7345 3991 7351 4017
rect 7377 3991 7383 4017
rect 6343 3985 6369 3991
rect 672 3933 9376 3950
rect 672 3907 2763 3933
rect 2789 3907 2815 3933
rect 2841 3907 2867 3933
rect 2893 3907 4919 3933
rect 4945 3907 4971 3933
rect 4997 3907 5023 3933
rect 5049 3907 7075 3933
rect 7101 3907 7127 3933
rect 7153 3907 7179 3933
rect 7205 3907 9231 3933
rect 9257 3907 9283 3933
rect 9309 3907 9335 3933
rect 9361 3907 9376 3933
rect 672 3890 9376 3907
rect 1807 3849 1833 3855
rect 7407 3849 7433 3855
rect 3985 3823 3991 3849
rect 4017 3823 4023 3849
rect 1807 3817 1833 3823
rect 7407 3817 7433 3823
rect 8135 3849 8161 3855
rect 8135 3817 8161 3823
rect 8751 3849 8777 3855
rect 8751 3817 8777 3823
rect 8863 3849 8889 3855
rect 8863 3817 8889 3823
rect 1023 3793 1049 3799
rect 1023 3761 1049 3767
rect 2479 3793 2505 3799
rect 2479 3761 2505 3767
rect 3375 3793 3401 3799
rect 8359 3793 8385 3799
rect 5441 3767 5447 3793
rect 5473 3767 5479 3793
rect 3375 3761 3401 3767
rect 8359 3761 8385 3767
rect 8975 3793 9001 3799
rect 8975 3761 9001 3767
rect 9031 3793 9057 3799
rect 9031 3761 9057 3767
rect 1079 3737 1105 3743
rect 1079 3705 1105 3711
rect 1527 3737 1553 3743
rect 1527 3705 1553 3711
rect 1751 3737 1777 3743
rect 1751 3705 1777 3711
rect 1863 3737 1889 3743
rect 1863 3705 1889 3711
rect 2031 3737 2057 3743
rect 2031 3705 2057 3711
rect 2199 3737 2225 3743
rect 2199 3705 2225 3711
rect 2311 3737 2337 3743
rect 3151 3737 3177 3743
rect 3033 3711 3039 3737
rect 3065 3711 3071 3737
rect 2311 3705 2337 3711
rect 3151 3705 3177 3711
rect 3543 3737 3569 3743
rect 8023 3737 8049 3743
rect 5497 3711 5503 3737
rect 5529 3711 5535 3737
rect 6169 3711 6175 3737
rect 6201 3711 6207 3737
rect 6953 3711 6959 3737
rect 6985 3711 6991 3737
rect 3543 3705 3569 3711
rect 8023 3705 8049 3711
rect 8247 3737 8273 3743
rect 8247 3705 8273 3711
rect 8695 3737 8721 3743
rect 8695 3705 8721 3711
rect 9143 3737 9169 3743
rect 9143 3705 9169 3711
rect 1247 3681 1273 3687
rect 1247 3649 1273 3655
rect 2255 3681 2281 3687
rect 2255 3649 2281 3655
rect 3711 3681 3737 3687
rect 6001 3655 6007 3681
rect 6033 3655 6039 3681
rect 3711 3649 3737 3655
rect 3207 3625 3233 3631
rect 3207 3593 3233 3599
rect 3823 3625 3849 3631
rect 3823 3593 3849 3599
rect 7295 3625 7321 3631
rect 7295 3593 7321 3599
rect 7463 3625 7489 3631
rect 7463 3593 7489 3599
rect 672 3541 9296 3558
rect 672 3515 1685 3541
rect 1711 3515 1737 3541
rect 1763 3515 1789 3541
rect 1815 3515 3841 3541
rect 3867 3515 3893 3541
rect 3919 3515 3945 3541
rect 3971 3515 5997 3541
rect 6023 3515 6049 3541
rect 6075 3515 6101 3541
rect 6127 3515 8153 3541
rect 8179 3515 8205 3541
rect 8231 3515 8257 3541
rect 8283 3515 9296 3541
rect 672 3498 9296 3515
rect 1415 3457 1441 3463
rect 3095 3457 3121 3463
rect 1577 3431 1583 3457
rect 1609 3431 1615 3457
rect 1415 3425 1441 3431
rect 3095 3425 3121 3431
rect 6287 3457 6313 3463
rect 6287 3425 6313 3431
rect 6455 3457 6481 3463
rect 7065 3431 7071 3457
rect 7097 3431 7103 3457
rect 6455 3425 6481 3431
rect 1303 3401 1329 3407
rect 1303 3369 1329 3375
rect 4271 3401 4297 3407
rect 6057 3375 6063 3401
rect 6089 3375 6095 3401
rect 6785 3375 6791 3401
rect 6817 3375 6823 3401
rect 9081 3375 9087 3401
rect 9113 3375 9119 3401
rect 4271 3369 4297 3375
rect 4047 3345 4073 3351
rect 2977 3319 2983 3345
rect 3009 3319 3015 3345
rect 3425 3319 3431 3345
rect 3457 3319 3463 3345
rect 3649 3319 3655 3345
rect 3681 3319 3687 3345
rect 4377 3319 4383 3345
rect 4409 3319 4415 3345
rect 4601 3319 4607 3345
rect 4633 3319 4639 3345
rect 6897 3319 6903 3345
rect 6929 3319 6935 3345
rect 7345 3319 7351 3345
rect 7377 3319 7383 3345
rect 7681 3319 7687 3345
rect 7713 3319 7719 3345
rect 8017 3319 8023 3345
rect 8049 3319 8055 3345
rect 4047 3313 4073 3319
rect 4153 3263 4159 3289
rect 4185 3263 4191 3289
rect 4993 3263 4999 3289
rect 5025 3263 5031 3289
rect 7457 3263 7463 3289
rect 7489 3263 7495 3289
rect 6399 3233 6425 3239
rect 4209 3207 4215 3233
rect 4241 3207 4247 3233
rect 6399 3201 6425 3207
rect 672 3149 9376 3166
rect 672 3123 2763 3149
rect 2789 3123 2815 3149
rect 2841 3123 2867 3149
rect 2893 3123 4919 3149
rect 4945 3123 4971 3149
rect 4997 3123 5023 3149
rect 5049 3123 7075 3149
rect 7101 3123 7127 3149
rect 7153 3123 7179 3149
rect 7205 3123 9231 3149
rect 9257 3123 9283 3149
rect 9309 3123 9335 3149
rect 9361 3123 9376 3149
rect 672 3106 9376 3123
rect 2815 3065 2841 3071
rect 2815 3033 2841 3039
rect 3095 3065 3121 3071
rect 3095 3033 3121 3039
rect 3207 3065 3233 3071
rect 3207 3033 3233 3039
rect 3487 3065 3513 3071
rect 3487 3033 3513 3039
rect 4439 3065 4465 3071
rect 4439 3033 4465 3039
rect 5223 3065 5249 3071
rect 5223 3033 5249 3039
rect 7911 3065 7937 3071
rect 7911 3033 7937 3039
rect 4999 3009 5025 3015
rect 1521 2983 1527 3009
rect 1553 2983 1559 3009
rect 4999 2977 5025 2983
rect 5279 3009 5305 3015
rect 6561 2983 6567 3009
rect 6593 2983 6599 3009
rect 5279 2977 5305 2983
rect 3039 2953 3065 2959
rect 3935 2953 3961 2959
rect 8639 2953 8665 2959
rect 1129 2927 1135 2953
rect 1161 2927 1167 2953
rect 3313 2927 3319 2953
rect 3345 2927 3351 2953
rect 3817 2927 3823 2953
rect 3849 2927 3855 2953
rect 6953 2927 6959 2953
rect 6985 2927 6991 2953
rect 8353 2927 8359 2953
rect 8385 2927 8391 2953
rect 3039 2921 3065 2927
rect 3935 2921 3961 2927
rect 8639 2921 8665 2927
rect 8863 2953 8889 2959
rect 8863 2921 8889 2927
rect 8919 2953 8945 2959
rect 8919 2921 8945 2927
rect 3151 2897 3177 2903
rect 8751 2897 8777 2903
rect 2585 2871 2591 2897
rect 2617 2871 2623 2897
rect 3873 2871 3879 2897
rect 3905 2871 3911 2897
rect 4993 2871 4999 2897
rect 5025 2871 5031 2897
rect 5497 2871 5503 2897
rect 5529 2871 5535 2897
rect 3151 2865 3177 2871
rect 8751 2865 8777 2871
rect 4887 2841 4913 2847
rect 4887 2809 4913 2815
rect 672 2757 9296 2774
rect 672 2731 1685 2757
rect 1711 2731 1737 2757
rect 1763 2731 1789 2757
rect 1815 2731 3841 2757
rect 3867 2731 3893 2757
rect 3919 2731 3945 2757
rect 3971 2731 5997 2757
rect 6023 2731 6049 2757
rect 6075 2731 6101 2757
rect 6127 2731 8153 2757
rect 8179 2731 8205 2757
rect 8231 2731 8257 2757
rect 8283 2731 9296 2757
rect 672 2714 9296 2731
rect 3095 2673 3121 2679
rect 3095 2641 3121 2647
rect 6959 2617 6985 2623
rect 9087 2617 9113 2623
rect 2921 2591 2927 2617
rect 2953 2591 2959 2617
rect 4937 2591 4943 2617
rect 4969 2591 4975 2617
rect 6001 2591 6007 2617
rect 6033 2591 6039 2617
rect 8465 2591 8471 2617
rect 8497 2591 8503 2617
rect 6959 2585 6985 2591
rect 9087 2585 9113 2591
rect 2591 2561 2617 2567
rect 2591 2529 2617 2535
rect 3431 2561 3457 2567
rect 6903 2561 6929 2567
rect 4097 2535 4103 2561
rect 4129 2535 4135 2561
rect 4321 2535 4327 2561
rect 4353 2535 4359 2561
rect 4769 2535 4775 2561
rect 4801 2535 4807 2561
rect 6393 2535 6399 2561
rect 6425 2535 6431 2561
rect 3431 2529 3457 2535
rect 6903 2529 6929 2535
rect 7015 2561 7041 2567
rect 7121 2535 7127 2561
rect 7153 2535 7159 2561
rect 8801 2535 8807 2561
rect 8833 2535 8839 2561
rect 7015 2529 7041 2535
rect 2983 2505 3009 2511
rect 3257 2479 3263 2505
rect 3289 2479 3295 2505
rect 2983 2473 3009 2479
rect 4719 2449 4745 2455
rect 4719 2417 4745 2423
rect 6847 2449 6873 2455
rect 7345 2423 7351 2449
rect 7377 2423 7383 2449
rect 6847 2417 6873 2423
rect 672 2365 9376 2382
rect 672 2339 2763 2365
rect 2789 2339 2815 2365
rect 2841 2339 2867 2365
rect 2893 2339 4919 2365
rect 4945 2339 4971 2365
rect 4997 2339 5023 2365
rect 5049 2339 7075 2365
rect 7101 2339 7127 2365
rect 7153 2339 7179 2365
rect 7205 2339 9231 2365
rect 9257 2339 9283 2365
rect 9309 2339 9335 2365
rect 9361 2339 9376 2365
rect 672 2322 9376 2339
rect 5111 2281 5137 2287
rect 5111 2249 5137 2255
rect 5223 2281 5249 2287
rect 6225 2255 6231 2281
rect 6257 2255 6263 2281
rect 5223 2249 5249 2255
rect 3991 2225 4017 2231
rect 2473 2199 2479 2225
rect 2505 2199 2511 2225
rect 3991 2193 4017 2199
rect 5447 2225 5473 2231
rect 6959 2225 6985 2231
rect 5609 2199 5615 2225
rect 5641 2199 5647 2225
rect 5447 2193 5473 2199
rect 6959 2193 6985 2199
rect 3823 2169 3849 2175
rect 2137 2143 2143 2169
rect 2169 2143 2175 2169
rect 3823 2137 3849 2143
rect 3935 2169 3961 2175
rect 3935 2137 3961 2143
rect 5279 2169 5305 2175
rect 5279 2137 5305 2143
rect 6343 2169 6369 2175
rect 8751 2169 8777 2175
rect 7233 2143 7239 2169
rect 7265 2143 7271 2169
rect 6343 2137 6369 2143
rect 8751 2137 8777 2143
rect 8695 2113 8721 2119
rect 3537 2087 3543 2113
rect 3569 2087 3575 2113
rect 8695 2081 8721 2087
rect 3767 2057 3793 2063
rect 3767 2025 3793 2031
rect 672 1973 9296 1990
rect 672 1947 1685 1973
rect 1711 1947 1737 1973
rect 1763 1947 1789 1973
rect 1815 1947 3841 1973
rect 3867 1947 3893 1973
rect 3919 1947 3945 1973
rect 3971 1947 5997 1973
rect 6023 1947 6049 1973
rect 6075 1947 6101 1973
rect 6127 1947 8153 1973
rect 8179 1947 8205 1973
rect 8231 1947 8257 1973
rect 8283 1947 9296 1973
rect 672 1930 9296 1947
rect 6623 1889 6649 1895
rect 6623 1857 6649 1863
rect 8079 1889 8105 1895
rect 8079 1857 8105 1863
rect 967 1833 993 1839
rect 967 1801 993 1807
rect 3711 1833 3737 1839
rect 3711 1801 3737 1807
rect 6175 1833 6201 1839
rect 6175 1801 6201 1807
rect 6679 1777 6705 1783
rect 1913 1751 1919 1777
rect 1945 1751 1951 1777
rect 5049 1751 5055 1777
rect 5081 1751 5087 1777
rect 7009 1751 7015 1777
rect 7041 1751 7047 1777
rect 6679 1745 6705 1751
rect 6623 1721 6649 1727
rect 6623 1689 6649 1695
rect 8807 1721 8833 1727
rect 8807 1689 8833 1695
rect 8919 1721 8945 1727
rect 8919 1689 8945 1695
rect 9087 1721 9113 1727
rect 9087 1689 9113 1695
rect 672 1581 9376 1598
rect 672 1555 2763 1581
rect 2789 1555 2815 1581
rect 2841 1555 2867 1581
rect 2893 1555 4919 1581
rect 4945 1555 4971 1581
rect 4997 1555 5023 1581
rect 5049 1555 7075 1581
rect 7101 1555 7127 1581
rect 7153 1555 7179 1581
rect 7205 1555 9231 1581
rect 9257 1555 9283 1581
rect 9309 1555 9335 1581
rect 9361 1555 9376 1581
rect 672 1538 9376 1555
<< via1 >>
rect 1685 8219 1711 8245
rect 1737 8219 1763 8245
rect 1789 8219 1815 8245
rect 3841 8219 3867 8245
rect 3893 8219 3919 8245
rect 3945 8219 3971 8245
rect 5997 8219 6023 8245
rect 6049 8219 6075 8245
rect 6101 8219 6127 8245
rect 8153 8219 8179 8245
rect 8205 8219 8231 8245
rect 8257 8219 8283 8245
rect 1247 8079 1273 8105
rect 8863 8079 8889 8105
rect 855 8023 881 8049
rect 8191 8023 8217 8049
rect 8583 8023 8609 8049
rect 6119 7967 6145 7993
rect 7407 7967 7433 7993
rect 1023 7911 1049 7937
rect 6287 7911 6313 7937
rect 8471 7911 8497 7937
rect 2763 7827 2789 7853
rect 2815 7827 2841 7853
rect 2867 7827 2893 7853
rect 4919 7827 4945 7853
rect 4971 7827 4997 7853
rect 5023 7827 5049 7853
rect 7075 7827 7101 7853
rect 7127 7827 7153 7853
rect 7179 7827 7205 7853
rect 9231 7827 9257 7853
rect 9283 7827 9309 7853
rect 9335 7827 9361 7853
rect 7911 7743 7937 7769
rect 8807 7743 8833 7769
rect 3039 7631 3065 7657
rect 3431 7631 3457 7657
rect 6903 7631 6929 7657
rect 8415 7631 8441 7657
rect 4495 7575 4521 7601
rect 4887 7575 4913 7601
rect 5447 7575 5473 7601
rect 6511 7575 6537 7601
rect 8807 7575 8833 7601
rect 8695 7519 8721 7545
rect 1685 7435 1711 7461
rect 1737 7435 1763 7461
rect 1789 7435 1815 7461
rect 3841 7435 3867 7461
rect 3893 7435 3919 7461
rect 3945 7435 3971 7461
rect 5997 7435 6023 7461
rect 6049 7435 6075 7461
rect 6101 7435 6127 7461
rect 8153 7435 8179 7461
rect 8205 7435 8231 7461
rect 8257 7435 8283 7461
rect 5951 7351 5977 7377
rect 4327 7295 4353 7321
rect 6399 7295 6425 7321
rect 9031 7295 9057 7321
rect 4551 7239 4577 7265
rect 4943 7239 4969 7265
rect 5111 7239 5137 7265
rect 5335 7239 5361 7265
rect 5895 7239 5921 7265
rect 7239 7239 7265 7265
rect 7295 7239 7321 7265
rect 7575 7239 7601 7265
rect 4775 7183 4801 7209
rect 4887 7183 4913 7209
rect 5559 7183 5585 7209
rect 6231 7183 6257 7209
rect 6455 7183 6481 7209
rect 7015 7183 7041 7209
rect 7127 7183 7153 7209
rect 7967 7183 7993 7209
rect 3935 7127 3961 7153
rect 4103 7127 4129 7153
rect 4439 7127 4465 7153
rect 5167 7127 5193 7153
rect 5615 7127 5641 7153
rect 5671 7127 5697 7153
rect 5727 7127 5753 7153
rect 6007 7127 6033 7153
rect 6119 7127 6145 7153
rect 7407 7127 7433 7153
rect 2763 7043 2789 7069
rect 2815 7043 2841 7069
rect 2867 7043 2893 7069
rect 4919 7043 4945 7069
rect 4971 7043 4997 7069
rect 5023 7043 5049 7069
rect 7075 7043 7101 7069
rect 7127 7043 7153 7069
rect 7179 7043 7205 7069
rect 9231 7043 9257 7069
rect 9283 7043 9309 7069
rect 9335 7043 9361 7069
rect 4551 6959 4577 6985
rect 6063 6959 6089 6985
rect 6679 6959 6705 6985
rect 6903 6959 6929 6985
rect 8751 6959 8777 6985
rect 4495 6903 4521 6929
rect 4775 6903 4801 6929
rect 2647 6847 2673 6873
rect 4271 6847 4297 6873
rect 4383 6847 4409 6873
rect 4887 6847 4913 6873
rect 4999 6847 5025 6873
rect 5839 6847 5865 6873
rect 5951 6847 5977 6873
rect 6175 6847 6201 6873
rect 6287 6847 6313 6873
rect 6399 6847 6425 6873
rect 6567 6847 6593 6873
rect 6959 6847 6985 6873
rect 8415 6847 8441 6873
rect 8863 6847 8889 6873
rect 2983 6791 3009 6817
rect 4047 6791 4073 6817
rect 6511 6791 6537 6817
rect 5111 6735 5137 6761
rect 5335 6735 5361 6761
rect 6063 6735 6089 6761
rect 6903 6735 6929 6761
rect 7911 6735 7937 6761
rect 8695 6735 8721 6761
rect 1685 6651 1711 6677
rect 1737 6651 1763 6677
rect 1789 6651 1815 6677
rect 3841 6651 3867 6677
rect 3893 6651 3919 6677
rect 3945 6651 3971 6677
rect 5997 6651 6023 6677
rect 6049 6651 6075 6677
rect 6101 6651 6127 6677
rect 8153 6651 8179 6677
rect 8205 6651 8231 6677
rect 8257 6651 8283 6677
rect 5055 6567 5081 6593
rect 5167 6567 5193 6593
rect 5783 6567 5809 6593
rect 4047 6511 4073 6537
rect 5335 6511 5361 6537
rect 8023 6511 8049 6537
rect 9087 6511 9113 6537
rect 4215 6455 4241 6481
rect 4719 6455 4745 6481
rect 5279 6455 5305 6481
rect 5671 6455 5697 6481
rect 5895 6455 5921 6481
rect 6007 6455 6033 6481
rect 7015 6455 7041 6481
rect 7631 6455 7657 6481
rect 855 6399 881 6425
rect 4439 6399 4465 6425
rect 4607 6399 4633 6425
rect 5559 6399 5585 6425
rect 6175 6399 6201 6425
rect 6343 6399 6369 6425
rect 7295 6399 7321 6425
rect 1023 6343 1049 6369
rect 1247 6343 1273 6369
rect 5335 6343 5361 6369
rect 5783 6343 5809 6369
rect 7127 6343 7153 6369
rect 7463 6343 7489 6369
rect 2763 6259 2789 6285
rect 2815 6259 2841 6285
rect 2867 6259 2893 6285
rect 4919 6259 4945 6285
rect 4971 6259 4997 6285
rect 5023 6259 5049 6285
rect 7075 6259 7101 6285
rect 7127 6259 7153 6285
rect 7179 6259 7205 6285
rect 9231 6259 9257 6285
rect 9283 6259 9309 6285
rect 9335 6259 9361 6285
rect 3599 6175 3625 6201
rect 3823 6175 3849 6201
rect 4047 6175 4073 6201
rect 4831 6175 4857 6201
rect 5223 6175 5249 6201
rect 4271 6119 4297 6145
rect 4495 6119 4521 6145
rect 5727 6119 5753 6145
rect 5951 6119 5977 6145
rect 6791 6119 6817 6145
rect 6959 6119 6985 6145
rect 1975 6063 2001 6089
rect 3991 6063 4017 6089
rect 4383 6063 4409 6089
rect 4999 6063 5025 6089
rect 5167 6063 5193 6089
rect 5335 6063 5361 6089
rect 5559 6063 5585 6089
rect 6399 6063 6425 6089
rect 8359 6063 8385 6089
rect 8639 6063 8665 6089
rect 8863 6063 8889 6089
rect 8919 6063 8945 6089
rect 2311 6007 2337 6033
rect 3375 6007 3401 6033
rect 6287 6007 6313 6033
rect 8751 6007 8777 6033
rect 4047 5951 4073 5977
rect 4551 5951 4577 5977
rect 5279 5951 5305 5977
rect 5895 5951 5921 5977
rect 6063 5951 6089 5977
rect 6231 5951 6257 5977
rect 7911 5951 7937 5977
rect 1685 5867 1711 5893
rect 1737 5867 1763 5893
rect 1789 5867 1815 5893
rect 3841 5867 3867 5893
rect 3893 5867 3919 5893
rect 3945 5867 3971 5893
rect 5997 5867 6023 5893
rect 6049 5867 6075 5893
rect 6101 5867 6127 5893
rect 8153 5867 8179 5893
rect 8205 5867 8231 5893
rect 8257 5867 8283 5893
rect 5167 5783 5193 5809
rect 5727 5783 5753 5809
rect 1415 5727 1441 5753
rect 1695 5727 1721 5753
rect 4271 5727 4297 5753
rect 4943 5727 4969 5753
rect 7295 5727 7321 5753
rect 8023 5727 8049 5753
rect 9087 5727 9113 5753
rect 1471 5671 1497 5697
rect 2815 5671 2841 5697
rect 4607 5671 4633 5697
rect 4887 5671 4913 5697
rect 4999 5671 5025 5697
rect 5167 5671 5193 5697
rect 6063 5671 6089 5697
rect 6343 5671 6369 5697
rect 6847 5671 6873 5697
rect 7183 5671 7209 5697
rect 7351 5671 7377 5697
rect 7631 5671 7657 5697
rect 3207 5615 3233 5641
rect 5895 5615 5921 5641
rect 6735 5615 6761 5641
rect 7071 5615 7097 5641
rect 1639 5559 1665 5585
rect 4439 5559 4465 5585
rect 5615 5559 5641 5585
rect 5671 5559 5697 5585
rect 6231 5559 6257 5585
rect 7463 5559 7489 5585
rect 2763 5475 2789 5501
rect 2815 5475 2841 5501
rect 2867 5475 2893 5501
rect 4919 5475 4945 5501
rect 4971 5475 4997 5501
rect 5023 5475 5049 5501
rect 7075 5475 7101 5501
rect 7127 5475 7153 5501
rect 7179 5475 7205 5501
rect 9231 5475 9257 5501
rect 9283 5475 9309 5501
rect 9335 5475 9361 5501
rect 1471 5391 1497 5417
rect 2535 5391 2561 5417
rect 2815 5391 2841 5417
rect 3151 5391 3177 5417
rect 7911 5391 7937 5417
rect 8751 5391 8777 5417
rect 8863 5391 8889 5417
rect 1415 5335 1441 5361
rect 2759 5335 2785 5361
rect 4271 5335 4297 5361
rect 4775 5335 4801 5361
rect 4831 5335 4857 5361
rect 7855 5335 7881 5361
rect 8191 5335 8217 5361
rect 1303 5279 1329 5305
rect 1639 5279 1665 5305
rect 2983 5279 3009 5305
rect 3207 5279 3233 5305
rect 3319 5279 3345 5305
rect 3487 5279 3513 5305
rect 3599 5279 3625 5305
rect 3767 5279 3793 5305
rect 3935 5279 3961 5305
rect 4495 5279 4521 5305
rect 4943 5279 4969 5305
rect 5111 5279 5137 5305
rect 8135 5279 8161 5305
rect 8303 5279 8329 5305
rect 8695 5279 8721 5305
rect 2871 5223 2897 5249
rect 3711 5223 3737 5249
rect 4439 5223 4465 5249
rect 6175 5223 6201 5249
rect 9031 5223 9057 5249
rect 1583 5167 1609 5193
rect 7911 5167 7937 5193
rect 1685 5083 1711 5109
rect 1737 5083 1763 5109
rect 1789 5083 1815 5109
rect 3841 5083 3867 5109
rect 3893 5083 3919 5109
rect 3945 5083 3971 5109
rect 5997 5083 6023 5109
rect 6049 5083 6075 5109
rect 6101 5083 6127 5109
rect 8153 5083 8179 5109
rect 8205 5083 8231 5109
rect 8257 5083 8283 5109
rect 6231 4999 6257 5025
rect 1471 4943 1497 4969
rect 2535 4943 2561 4969
rect 3655 4943 3681 4969
rect 8975 4943 9001 4969
rect 1135 4887 1161 4913
rect 5727 4887 5753 4913
rect 5951 4887 5977 4913
rect 6343 4887 6369 4913
rect 6847 4887 6873 4913
rect 7127 4887 7153 4913
rect 7575 4887 7601 4913
rect 6063 4831 6089 4857
rect 7295 4831 7321 4857
rect 7911 4831 7937 4857
rect 2983 4775 3009 4801
rect 6343 4775 6369 4801
rect 6959 4775 6985 4801
rect 2763 4691 2789 4717
rect 2815 4691 2841 4717
rect 2867 4691 2893 4717
rect 4919 4691 4945 4717
rect 4971 4691 4997 4717
rect 5023 4691 5049 4717
rect 7075 4691 7101 4717
rect 7127 4691 7153 4717
rect 7179 4691 7205 4717
rect 9231 4691 9257 4717
rect 9283 4691 9309 4717
rect 9335 4691 9361 4717
rect 2647 4607 2673 4633
rect 4831 4607 4857 4633
rect 8751 4607 8777 4633
rect 2759 4551 2785 4577
rect 3375 4551 3401 4577
rect 4775 4551 4801 4577
rect 5615 4551 5641 4577
rect 7575 4551 7601 4577
rect 8695 4551 8721 4577
rect 8975 4551 9001 4577
rect 1135 4495 1161 4521
rect 2815 4495 2841 4521
rect 3039 4495 3065 4521
rect 5335 4495 5361 4521
rect 5783 4495 5809 4521
rect 8863 4495 8889 4521
rect 911 4439 937 4465
rect 1471 4439 1497 4465
rect 2535 4439 2561 4465
rect 4439 4439 4465 4465
rect 5391 4439 5417 4465
rect 4831 4383 4857 4409
rect 1685 4299 1711 4325
rect 1737 4299 1763 4325
rect 1789 4299 1815 4325
rect 3841 4299 3867 4325
rect 3893 4299 3919 4325
rect 3945 4299 3971 4325
rect 5997 4299 6023 4325
rect 6049 4299 6075 4325
rect 6101 4299 6127 4325
rect 8153 4299 8179 4325
rect 8205 4299 8231 4325
rect 8257 4299 8283 4325
rect 1583 4215 1609 4241
rect 5951 4215 5977 4241
rect 1919 4159 1945 4185
rect 2871 4159 2897 4185
rect 3711 4159 3737 4185
rect 4551 4159 4577 4185
rect 6735 4159 6761 4185
rect 9087 4159 9113 4185
rect 911 4103 937 4129
rect 1415 4103 1441 4129
rect 1583 4103 1609 4129
rect 1975 4103 2001 4129
rect 2143 4103 2169 4129
rect 5223 4103 5249 4129
rect 5391 4103 5417 4129
rect 6847 4103 6873 4129
rect 7239 4103 7265 4129
rect 7687 4103 7713 4129
rect 1303 4047 1329 4073
rect 1863 4047 1889 4073
rect 4943 4047 4969 4073
rect 5895 4047 5921 4073
rect 6287 4047 6313 4073
rect 6399 4047 6425 4073
rect 8023 4047 8049 4073
rect 1023 3991 1049 4017
rect 1471 3991 1497 4017
rect 3655 3991 3681 4017
rect 3767 3991 3793 4017
rect 3879 3991 3905 4017
rect 6343 3991 6369 4017
rect 7015 3991 7041 4017
rect 7351 3991 7377 4017
rect 2763 3907 2789 3933
rect 2815 3907 2841 3933
rect 2867 3907 2893 3933
rect 4919 3907 4945 3933
rect 4971 3907 4997 3933
rect 5023 3907 5049 3933
rect 7075 3907 7101 3933
rect 7127 3907 7153 3933
rect 7179 3907 7205 3933
rect 9231 3907 9257 3933
rect 9283 3907 9309 3933
rect 9335 3907 9361 3933
rect 1807 3823 1833 3849
rect 3991 3823 4017 3849
rect 7407 3823 7433 3849
rect 8135 3823 8161 3849
rect 8751 3823 8777 3849
rect 8863 3823 8889 3849
rect 1023 3767 1049 3793
rect 2479 3767 2505 3793
rect 3375 3767 3401 3793
rect 5447 3767 5473 3793
rect 8359 3767 8385 3793
rect 8975 3767 9001 3793
rect 9031 3767 9057 3793
rect 1079 3711 1105 3737
rect 1527 3711 1553 3737
rect 1751 3711 1777 3737
rect 1863 3711 1889 3737
rect 2031 3711 2057 3737
rect 2199 3711 2225 3737
rect 2311 3711 2337 3737
rect 3039 3711 3065 3737
rect 3151 3711 3177 3737
rect 3543 3711 3569 3737
rect 5503 3711 5529 3737
rect 6175 3711 6201 3737
rect 6959 3711 6985 3737
rect 8023 3711 8049 3737
rect 8247 3711 8273 3737
rect 8695 3711 8721 3737
rect 9143 3711 9169 3737
rect 1247 3655 1273 3681
rect 2255 3655 2281 3681
rect 3711 3655 3737 3681
rect 6007 3655 6033 3681
rect 3207 3599 3233 3625
rect 3823 3599 3849 3625
rect 7295 3599 7321 3625
rect 7463 3599 7489 3625
rect 1685 3515 1711 3541
rect 1737 3515 1763 3541
rect 1789 3515 1815 3541
rect 3841 3515 3867 3541
rect 3893 3515 3919 3541
rect 3945 3515 3971 3541
rect 5997 3515 6023 3541
rect 6049 3515 6075 3541
rect 6101 3515 6127 3541
rect 8153 3515 8179 3541
rect 8205 3515 8231 3541
rect 8257 3515 8283 3541
rect 1415 3431 1441 3457
rect 1583 3431 1609 3457
rect 3095 3431 3121 3457
rect 6287 3431 6313 3457
rect 6455 3431 6481 3457
rect 7071 3431 7097 3457
rect 1303 3375 1329 3401
rect 4271 3375 4297 3401
rect 6063 3375 6089 3401
rect 6791 3375 6817 3401
rect 9087 3375 9113 3401
rect 2983 3319 3009 3345
rect 3431 3319 3457 3345
rect 3655 3319 3681 3345
rect 4047 3319 4073 3345
rect 4383 3319 4409 3345
rect 4607 3319 4633 3345
rect 6903 3319 6929 3345
rect 7351 3319 7377 3345
rect 7687 3319 7713 3345
rect 8023 3319 8049 3345
rect 4159 3263 4185 3289
rect 4999 3263 5025 3289
rect 7463 3263 7489 3289
rect 4215 3207 4241 3233
rect 6399 3207 6425 3233
rect 2763 3123 2789 3149
rect 2815 3123 2841 3149
rect 2867 3123 2893 3149
rect 4919 3123 4945 3149
rect 4971 3123 4997 3149
rect 5023 3123 5049 3149
rect 7075 3123 7101 3149
rect 7127 3123 7153 3149
rect 7179 3123 7205 3149
rect 9231 3123 9257 3149
rect 9283 3123 9309 3149
rect 9335 3123 9361 3149
rect 2815 3039 2841 3065
rect 3095 3039 3121 3065
rect 3207 3039 3233 3065
rect 3487 3039 3513 3065
rect 4439 3039 4465 3065
rect 5223 3039 5249 3065
rect 7911 3039 7937 3065
rect 1527 2983 1553 3009
rect 4999 2983 5025 3009
rect 5279 2983 5305 3009
rect 6567 2983 6593 3009
rect 1135 2927 1161 2953
rect 3039 2927 3065 2953
rect 3319 2927 3345 2953
rect 3823 2927 3849 2953
rect 3935 2927 3961 2953
rect 6959 2927 6985 2953
rect 8359 2927 8385 2953
rect 8639 2927 8665 2953
rect 8863 2927 8889 2953
rect 8919 2927 8945 2953
rect 2591 2871 2617 2897
rect 3151 2871 3177 2897
rect 3879 2871 3905 2897
rect 4999 2871 5025 2897
rect 5503 2871 5529 2897
rect 8751 2871 8777 2897
rect 4887 2815 4913 2841
rect 1685 2731 1711 2757
rect 1737 2731 1763 2757
rect 1789 2731 1815 2757
rect 3841 2731 3867 2757
rect 3893 2731 3919 2757
rect 3945 2731 3971 2757
rect 5997 2731 6023 2757
rect 6049 2731 6075 2757
rect 6101 2731 6127 2757
rect 8153 2731 8179 2757
rect 8205 2731 8231 2757
rect 8257 2731 8283 2757
rect 3095 2647 3121 2673
rect 2927 2591 2953 2617
rect 4943 2591 4969 2617
rect 6007 2591 6033 2617
rect 6959 2591 6985 2617
rect 8471 2591 8497 2617
rect 9087 2591 9113 2617
rect 2591 2535 2617 2561
rect 3431 2535 3457 2561
rect 4103 2535 4129 2561
rect 4327 2535 4353 2561
rect 4775 2535 4801 2561
rect 6399 2535 6425 2561
rect 6903 2535 6929 2561
rect 7015 2535 7041 2561
rect 7127 2535 7153 2561
rect 8807 2535 8833 2561
rect 2983 2479 3009 2505
rect 3263 2479 3289 2505
rect 4719 2423 4745 2449
rect 6847 2423 6873 2449
rect 7351 2423 7377 2449
rect 2763 2339 2789 2365
rect 2815 2339 2841 2365
rect 2867 2339 2893 2365
rect 4919 2339 4945 2365
rect 4971 2339 4997 2365
rect 5023 2339 5049 2365
rect 7075 2339 7101 2365
rect 7127 2339 7153 2365
rect 7179 2339 7205 2365
rect 9231 2339 9257 2365
rect 9283 2339 9309 2365
rect 9335 2339 9361 2365
rect 5111 2255 5137 2281
rect 5223 2255 5249 2281
rect 6231 2255 6257 2281
rect 2479 2199 2505 2225
rect 3991 2199 4017 2225
rect 5447 2199 5473 2225
rect 5615 2199 5641 2225
rect 6959 2199 6985 2225
rect 2143 2143 2169 2169
rect 3823 2143 3849 2169
rect 3935 2143 3961 2169
rect 5279 2143 5305 2169
rect 6343 2143 6369 2169
rect 7239 2143 7265 2169
rect 8751 2143 8777 2169
rect 3543 2087 3569 2113
rect 8695 2087 8721 2113
rect 3767 2031 3793 2057
rect 1685 1947 1711 1973
rect 1737 1947 1763 1973
rect 1789 1947 1815 1973
rect 3841 1947 3867 1973
rect 3893 1947 3919 1973
rect 3945 1947 3971 1973
rect 5997 1947 6023 1973
rect 6049 1947 6075 1973
rect 6101 1947 6127 1973
rect 8153 1947 8179 1973
rect 8205 1947 8231 1973
rect 8257 1947 8283 1973
rect 6623 1863 6649 1889
rect 8079 1863 8105 1889
rect 967 1807 993 1833
rect 3711 1807 3737 1833
rect 6175 1807 6201 1833
rect 1919 1751 1945 1777
rect 5055 1751 5081 1777
rect 6679 1751 6705 1777
rect 7015 1751 7041 1777
rect 6623 1695 6649 1721
rect 8807 1695 8833 1721
rect 8919 1695 8945 1721
rect 9087 1695 9113 1721
rect 2763 1555 2789 1581
rect 2815 1555 2841 1581
rect 2867 1555 2893 1581
rect 4919 1555 4945 1581
rect 4971 1555 4997 1581
rect 5023 1555 5049 1581
rect 7075 1555 7101 1581
rect 7127 1555 7153 1581
rect 7179 1555 7205 1581
rect 9231 1555 9257 1581
rect 9283 1555 9309 1581
rect 9335 1555 9361 1581
<< metal2 >>
rect 2464 9600 2520 10000
rect 7392 9600 7448 10000
rect 854 8666 882 8671
rect 854 8106 882 8638
rect 1684 8246 1816 8251
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1684 8213 1816 8218
rect 854 8049 882 8078
rect 1246 8106 1274 8111
rect 1246 8059 1274 8078
rect 854 8023 855 8049
rect 881 8023 882 8049
rect 854 8017 882 8023
rect 1022 7938 1050 7943
rect 1022 7891 1050 7910
rect 1862 7938 1890 7943
rect 1684 7462 1816 7467
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1684 7429 1816 7434
rect 1684 6678 1816 6683
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1684 6645 1816 6650
rect 854 6425 882 6431
rect 854 6399 855 6425
rect 881 6399 882 6425
rect 854 6202 882 6399
rect 1022 6370 1050 6375
rect 1022 6369 1218 6370
rect 1022 6343 1023 6369
rect 1049 6343 1218 6369
rect 1022 6342 1218 6343
rect 1022 6337 1050 6342
rect 854 6169 882 6174
rect 1190 5978 1218 6342
rect 1246 6369 1274 6375
rect 1246 6343 1247 6369
rect 1273 6343 1274 6369
rect 1246 6202 1274 6343
rect 1246 6169 1274 6174
rect 1190 5950 1442 5978
rect 1414 5753 1442 5950
rect 1684 5894 1816 5899
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1684 5861 1816 5866
rect 1862 5810 1890 7910
rect 2478 6202 2506 9600
rect 7406 8386 7434 9600
rect 7406 8353 7434 8358
rect 7910 9226 7938 9231
rect 3840 8246 3972 8251
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3840 8213 3972 8218
rect 5996 8246 6128 8251
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 5996 8213 6128 8218
rect 5446 7994 5474 7999
rect 2762 7854 2894 7859
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2762 7821 2894 7826
rect 4918 7854 5050 7859
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 4918 7821 5050 7826
rect 3038 7658 3066 7663
rect 2926 7657 3066 7658
rect 2926 7631 3039 7657
rect 3065 7631 3066 7657
rect 2926 7630 3066 7631
rect 2926 7574 2954 7630
rect 3038 7625 3066 7630
rect 3430 7658 3458 7663
rect 3430 7611 3458 7630
rect 4494 7601 4522 7607
rect 4886 7602 4914 7607
rect 4494 7575 4495 7601
rect 4521 7575 4522 7601
rect 2646 7546 3122 7574
rect 2646 6874 2674 7546
rect 3094 7378 3122 7546
rect 4494 7490 4522 7575
rect 3840 7462 3972 7467
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 4494 7457 4522 7462
rect 4550 7601 4914 7602
rect 4550 7575 4887 7601
rect 4913 7575 4914 7601
rect 4550 7574 4914 7575
rect 3840 7429 3972 7434
rect 3094 7345 3122 7350
rect 3598 7378 3626 7383
rect 3374 7154 3402 7159
rect 2762 7070 2894 7075
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2762 7037 2894 7042
rect 2646 6873 2730 6874
rect 2646 6847 2647 6873
rect 2673 6847 2730 6873
rect 2646 6846 2730 6847
rect 2646 6841 2674 6846
rect 2478 6169 2506 6174
rect 1974 6090 2002 6095
rect 1974 6043 2002 6062
rect 2702 6090 2730 6846
rect 2982 6818 3010 6823
rect 2982 6771 3010 6790
rect 2762 6286 2894 6291
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2762 6253 2894 6258
rect 2310 6033 2338 6039
rect 2310 6007 2311 6033
rect 2337 6007 2338 6033
rect 2310 5978 2338 6007
rect 2310 5945 2338 5950
rect 1414 5727 1415 5753
rect 1441 5727 1442 5753
rect 1414 5721 1442 5727
rect 1694 5782 1890 5810
rect 1694 5753 1722 5782
rect 2702 5754 2730 6062
rect 3374 6033 3402 7126
rect 3598 6202 3626 7350
rect 4326 7378 4354 7383
rect 4550 7378 4578 7574
rect 4886 7569 4914 7574
rect 4942 7602 4970 7607
rect 4774 7490 4802 7495
rect 4354 7350 4578 7378
rect 4718 7462 4774 7490
rect 4326 7321 4354 7350
rect 4326 7295 4327 7321
rect 4353 7295 4354 7321
rect 4326 7289 4354 7295
rect 4550 7266 4578 7271
rect 4494 7265 4578 7266
rect 4494 7239 4551 7265
rect 4577 7239 4578 7265
rect 4494 7238 4578 7239
rect 3934 7154 3962 7159
rect 3934 7107 3962 7126
rect 4102 7153 4130 7159
rect 4102 7127 4103 7153
rect 4129 7127 4130 7153
rect 4046 6817 4074 6823
rect 4046 6791 4047 6817
rect 4073 6791 4074 6817
rect 4046 6762 4074 6791
rect 4102 6762 4130 7127
rect 4438 7153 4466 7159
rect 4438 7127 4439 7153
rect 4465 7127 4466 7153
rect 4438 7098 4466 7127
rect 4326 7070 4466 7098
rect 4270 6873 4298 6879
rect 4270 6847 4271 6873
rect 4297 6847 4298 6873
rect 4102 6734 4242 6762
rect 3840 6678 3972 6683
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3840 6645 3972 6650
rect 4046 6537 4074 6734
rect 4046 6511 4047 6537
rect 4073 6511 4074 6537
rect 4046 6505 4074 6511
rect 4214 6482 4242 6734
rect 4214 6435 4242 6454
rect 4046 6426 4074 6431
rect 3822 6202 3850 6207
rect 3598 6201 3850 6202
rect 3598 6175 3599 6201
rect 3625 6175 3823 6201
rect 3849 6175 3850 6201
rect 3598 6174 3850 6175
rect 3598 6169 3626 6174
rect 3374 6007 3375 6033
rect 3401 6007 3402 6033
rect 3374 6001 3402 6007
rect 1694 5727 1695 5753
rect 1721 5727 1722 5753
rect 1694 5721 1722 5727
rect 2534 5726 2842 5754
rect 1470 5697 1498 5703
rect 1470 5671 1471 5697
rect 1497 5671 1498 5697
rect 1470 5642 1498 5671
rect 1358 5614 1498 5642
rect 1302 5305 1330 5311
rect 1302 5279 1303 5305
rect 1329 5279 1330 5305
rect 1134 4913 1162 4919
rect 1134 4887 1135 4913
rect 1161 4887 1162 4913
rect 1134 4521 1162 4887
rect 1134 4495 1135 4521
rect 1161 4495 1162 4521
rect 910 4465 938 4471
rect 910 4439 911 4465
rect 937 4439 938 4465
rect 910 4129 938 4439
rect 910 4103 911 4129
rect 937 4103 938 4129
rect 910 3738 938 4103
rect 1022 4017 1050 4023
rect 1022 3991 1023 4017
rect 1049 3991 1050 4017
rect 1022 3794 1050 3991
rect 1022 3747 1050 3766
rect 910 3705 938 3710
rect 1078 3738 1106 3743
rect 1078 3691 1106 3710
rect 1134 2954 1162 4495
rect 1302 4074 1330 5279
rect 1358 4130 1386 5614
rect 1638 5586 1666 5591
rect 1414 5585 1666 5586
rect 1414 5559 1639 5585
rect 1665 5559 1666 5585
rect 1414 5558 1666 5559
rect 1414 5361 1442 5558
rect 1638 5553 1666 5558
rect 1638 5474 1666 5479
rect 1414 5335 1415 5361
rect 1441 5335 1442 5361
rect 1414 5329 1442 5335
rect 1470 5417 1498 5423
rect 1470 5391 1471 5417
rect 1497 5391 1498 5417
rect 1470 4969 1498 5391
rect 1638 5306 1666 5446
rect 2534 5417 2562 5726
rect 2814 5697 2842 5726
rect 2814 5671 2815 5697
rect 2841 5671 2842 5697
rect 2814 5665 2842 5671
rect 3206 5642 3234 5647
rect 2926 5641 3234 5642
rect 2926 5615 3207 5641
rect 3233 5615 3234 5641
rect 2926 5614 3234 5615
rect 2762 5502 2894 5507
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2762 5469 2894 5474
rect 2534 5391 2535 5417
rect 2561 5391 2562 5417
rect 2534 5385 2562 5391
rect 2814 5418 2842 5423
rect 2926 5418 2954 5614
rect 3206 5609 3234 5614
rect 2814 5417 2954 5418
rect 2814 5391 2815 5417
rect 2841 5391 2954 5417
rect 2814 5390 2954 5391
rect 3150 5418 3178 5423
rect 3318 5418 3346 5423
rect 3150 5417 3290 5418
rect 3150 5391 3151 5417
rect 3177 5391 3290 5417
rect 3150 5390 3290 5391
rect 2814 5385 2842 5390
rect 3150 5385 3178 5390
rect 2758 5361 2786 5367
rect 2758 5335 2759 5361
rect 2785 5335 2786 5361
rect 1470 4943 1471 4969
rect 1497 4943 1498 4969
rect 1470 4937 1498 4943
rect 1526 5305 1666 5306
rect 1526 5279 1639 5305
rect 1665 5279 1666 5305
rect 1526 5278 1666 5279
rect 1470 4465 1498 4471
rect 1470 4439 1471 4465
rect 1497 4439 1498 4465
rect 1414 4130 1442 4135
rect 1358 4129 1442 4130
rect 1358 4103 1415 4129
rect 1441 4103 1442 4129
rect 1358 4102 1442 4103
rect 1414 4097 1442 4102
rect 1246 4073 1330 4074
rect 1246 4047 1303 4073
rect 1329 4047 1330 4073
rect 1246 4046 1330 4047
rect 1246 3681 1274 4046
rect 1302 4041 1330 4046
rect 1470 4017 1498 4439
rect 1526 4130 1554 5278
rect 1638 5273 1666 5278
rect 2590 5306 2618 5311
rect 1582 5193 1610 5199
rect 1582 5167 1583 5193
rect 1609 5167 1610 5193
rect 1582 4746 1610 5167
rect 1684 5110 1816 5115
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1684 5077 1816 5082
rect 2534 4969 2562 4975
rect 2534 4943 2535 4969
rect 2561 4943 2562 4969
rect 1582 4718 1946 4746
rect 1684 4326 1816 4331
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1684 4293 1816 4298
rect 1582 4241 1610 4247
rect 1582 4215 1583 4241
rect 1609 4215 1610 4241
rect 1582 4214 1610 4215
rect 1582 4186 1834 4214
rect 1582 4130 1610 4135
rect 1526 4129 1610 4130
rect 1526 4103 1583 4129
rect 1609 4103 1610 4129
rect 1526 4102 1610 4103
rect 1582 4097 1610 4102
rect 1470 3991 1471 4017
rect 1497 3991 1498 4017
rect 1470 3985 1498 3991
rect 1750 4074 1778 4079
rect 1246 3655 1247 3681
rect 1273 3655 1274 3681
rect 1246 3290 1274 3655
rect 1302 3794 1330 3799
rect 1302 3401 1330 3766
rect 1526 3738 1554 3743
rect 1526 3737 1610 3738
rect 1526 3711 1527 3737
rect 1553 3711 1610 3737
rect 1526 3710 1610 3711
rect 1526 3705 1554 3710
rect 1414 3682 1442 3687
rect 1414 3457 1442 3654
rect 1414 3431 1415 3457
rect 1441 3431 1442 3457
rect 1414 3425 1442 3431
rect 1582 3457 1610 3710
rect 1750 3737 1778 4046
rect 1806 3849 1834 4186
rect 1918 4185 1946 4718
rect 1918 4159 1919 4185
rect 1945 4159 1946 4185
rect 1918 4153 1946 4159
rect 2142 4578 2170 4583
rect 1974 4129 2002 4135
rect 1974 4103 1975 4129
rect 2001 4103 2002 4129
rect 1862 4074 1890 4079
rect 1862 4027 1890 4046
rect 1806 3823 1807 3849
rect 1833 3823 1834 3849
rect 1806 3817 1834 3823
rect 1750 3711 1751 3737
rect 1777 3711 1778 3737
rect 1750 3682 1778 3711
rect 1862 3794 1890 3799
rect 1974 3794 2002 4103
rect 2142 4129 2170 4550
rect 2534 4578 2562 4943
rect 2534 4545 2562 4550
rect 2590 4522 2618 5278
rect 2702 5026 2730 5031
rect 2646 4998 2702 5026
rect 2646 4633 2674 4998
rect 2702 4993 2730 4998
rect 2758 4970 2786 5335
rect 2982 5305 3010 5311
rect 2982 5279 2983 5305
rect 3009 5279 3010 5305
rect 2870 5250 2898 5255
rect 2870 5203 2898 5222
rect 2982 5026 3010 5279
rect 3206 5305 3234 5311
rect 3206 5279 3207 5305
rect 3233 5279 3234 5305
rect 2982 4993 3010 4998
rect 3094 5082 3122 5087
rect 3038 4970 3066 4975
rect 2758 4942 2842 4970
rect 2814 4858 2842 4942
rect 2814 4830 3010 4858
rect 2982 4801 3010 4830
rect 2982 4775 2983 4801
rect 3009 4775 3010 4801
rect 2762 4718 2894 4723
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2762 4685 2894 4690
rect 2646 4607 2647 4633
rect 2673 4607 2674 4633
rect 2646 4601 2674 4607
rect 2758 4578 2786 4583
rect 2758 4531 2786 4550
rect 2590 4494 2730 4522
rect 2142 4103 2143 4129
rect 2169 4103 2170 4129
rect 2142 4097 2170 4103
rect 2534 4465 2562 4471
rect 2534 4439 2535 4465
rect 2561 4439 2562 4465
rect 1890 3766 2002 3794
rect 2478 3794 2506 3799
rect 1862 3737 1890 3766
rect 2478 3747 2506 3766
rect 1862 3711 1863 3737
rect 1889 3711 1890 3737
rect 1862 3705 1890 3711
rect 2030 3737 2058 3743
rect 2030 3711 2031 3737
rect 2057 3711 2058 3737
rect 1750 3649 1778 3654
rect 1684 3542 1816 3547
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1684 3509 1816 3514
rect 2030 3514 2058 3711
rect 2030 3481 2058 3486
rect 2198 3737 2226 3743
rect 2198 3711 2199 3737
rect 2225 3711 2226 3737
rect 2198 3682 2226 3711
rect 2310 3738 2338 3743
rect 2310 3691 2338 3710
rect 1582 3431 1583 3457
rect 1609 3431 1610 3457
rect 1582 3425 1610 3431
rect 2198 3458 2226 3654
rect 2198 3425 2226 3430
rect 2254 3681 2282 3687
rect 2254 3655 2255 3681
rect 2281 3655 2282 3681
rect 1302 3375 1303 3401
rect 1329 3375 1330 3401
rect 1302 3369 1330 3375
rect 1526 3402 1554 3407
rect 1302 3290 1330 3295
rect 1246 3262 1302 3290
rect 1302 3257 1330 3262
rect 1526 3009 1554 3374
rect 2254 3402 2282 3655
rect 2534 3514 2562 4439
rect 2534 3481 2562 3486
rect 2702 4466 2730 4494
rect 2814 4521 2842 4527
rect 2814 4495 2815 4521
rect 2841 4495 2842 4521
rect 2814 4466 2842 4495
rect 2702 4438 2842 4466
rect 2870 4522 2898 4527
rect 2254 3369 2282 3374
rect 1526 2983 1527 3009
rect 1553 2983 1554 3009
rect 1526 2977 1554 2983
rect 1918 3290 1946 3295
rect 1134 2907 1162 2926
rect 1684 2758 1816 2763
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1684 2725 1816 2730
rect 1684 1974 1816 1979
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1684 1941 1816 1946
rect 966 1833 994 1839
rect 966 1807 967 1833
rect 993 1807 994 1833
rect 966 1274 994 1807
rect 1918 1777 1946 3262
rect 2702 3066 2730 4438
rect 2870 4186 2898 4494
rect 2870 4185 2954 4186
rect 2870 4159 2871 4185
rect 2897 4159 2954 4185
rect 2870 4158 2954 4159
rect 2870 4153 2898 4158
rect 2762 3934 2894 3939
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2762 3901 2894 3906
rect 2762 3150 2894 3155
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2762 3117 2894 3122
rect 2702 3033 2730 3038
rect 2814 3066 2842 3071
rect 2926 3066 2954 4158
rect 2982 3850 3010 4775
rect 3038 4522 3066 4942
rect 3038 4475 3066 4494
rect 2982 3817 3010 3822
rect 3094 3794 3122 5054
rect 3206 4634 3234 5279
rect 3206 4601 3234 4606
rect 3262 4578 3290 5390
rect 3318 5305 3346 5390
rect 3318 5279 3319 5305
rect 3345 5279 3346 5305
rect 3318 5082 3346 5279
rect 3486 5306 3514 5311
rect 3486 5259 3514 5278
rect 3598 5306 3626 5311
rect 3598 5259 3626 5278
rect 3318 5049 3346 5054
rect 3654 4970 3682 6174
rect 3822 6169 3850 6174
rect 4046 6201 4074 6398
rect 4270 6426 4298 6847
rect 4270 6393 4298 6398
rect 4326 6314 4354 7070
rect 4494 7042 4522 7238
rect 4550 7233 4578 7238
rect 4662 7210 4690 7215
rect 4438 7014 4522 7042
rect 4606 7182 4662 7210
rect 4382 6873 4410 6879
rect 4382 6847 4383 6873
rect 4409 6847 4410 6873
rect 4382 6538 4410 6847
rect 4438 6762 4466 7014
rect 4550 6986 4578 6991
rect 4606 6986 4634 7182
rect 4662 7177 4690 7182
rect 4550 6985 4634 6986
rect 4550 6959 4551 6985
rect 4577 6959 4634 6985
rect 4550 6958 4634 6959
rect 4550 6953 4578 6958
rect 4494 6930 4522 6935
rect 4718 6930 4746 7462
rect 4774 7457 4802 7462
rect 4942 7378 4970 7574
rect 5446 7602 5474 7966
rect 6118 7994 6146 7999
rect 6118 7947 6146 7966
rect 7406 7994 7434 7999
rect 7406 7947 7434 7966
rect 6286 7938 6314 7943
rect 6286 7937 6426 7938
rect 6286 7911 6287 7937
rect 6313 7911 6426 7937
rect 6286 7910 6426 7911
rect 6286 7905 6314 7910
rect 5446 7555 5474 7574
rect 5782 7658 5810 7663
rect 4886 7350 4970 7378
rect 4998 7490 5026 7495
rect 4774 7209 4802 7215
rect 4886 7210 4914 7350
rect 4942 7266 4970 7271
rect 4998 7266 5026 7462
rect 5110 7266 5138 7271
rect 5278 7266 5306 7271
rect 4942 7265 5138 7266
rect 4942 7239 4943 7265
rect 4969 7239 5111 7265
rect 5137 7239 5138 7265
rect 4942 7238 5138 7239
rect 4942 7233 4970 7238
rect 4774 7183 4775 7209
rect 4801 7183 4802 7209
rect 4774 7154 4802 7183
rect 4774 7121 4802 7126
rect 4830 7209 4914 7210
rect 4830 7183 4887 7209
rect 4913 7183 4914 7209
rect 4830 7182 4914 7183
rect 4774 6930 4802 6935
rect 4718 6929 4802 6930
rect 4718 6903 4775 6929
rect 4801 6903 4802 6929
rect 4718 6902 4802 6903
rect 4494 6883 4522 6902
rect 4774 6897 4802 6902
rect 4830 6874 4858 7182
rect 4886 7177 4914 7182
rect 4918 7070 5050 7075
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 4918 7037 5050 7042
rect 4998 6986 5026 6991
rect 5110 6986 5138 7238
rect 5222 7238 5278 7266
rect 5166 7154 5194 7159
rect 5166 7107 5194 7126
rect 5222 7042 5250 7238
rect 5278 7233 5306 7238
rect 5334 7265 5362 7271
rect 5334 7239 5335 7265
rect 5361 7239 5362 7265
rect 4886 6874 4914 6879
rect 4830 6873 4914 6874
rect 4830 6847 4887 6873
rect 4913 6847 4914 6873
rect 4830 6846 4914 6847
rect 4886 6841 4914 6846
rect 4998 6873 5026 6958
rect 4998 6847 4999 6873
rect 5025 6847 5026 6873
rect 4998 6841 5026 6847
rect 5054 6958 5138 6986
rect 5166 7014 5250 7042
rect 4438 6729 4466 6734
rect 4718 6762 4746 6767
rect 4662 6594 4690 6599
rect 4382 6505 4410 6510
rect 4606 6538 4634 6543
rect 4438 6426 4466 6431
rect 4046 6175 4047 6201
rect 4073 6175 4074 6201
rect 4046 6169 4074 6175
rect 4214 6286 4354 6314
rect 4382 6425 4466 6426
rect 4382 6399 4439 6425
rect 4465 6399 4466 6425
rect 4382 6398 4466 6399
rect 3990 6090 4018 6095
rect 3990 6043 4018 6062
rect 4046 5977 4074 5983
rect 4046 5951 4047 5977
rect 4073 5951 4074 5977
rect 3840 5894 3972 5899
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3840 5861 3972 5866
rect 3766 5305 3794 5311
rect 3766 5279 3767 5305
rect 3793 5279 3794 5305
rect 3710 5250 3738 5255
rect 3710 5203 3738 5222
rect 3654 4923 3682 4942
rect 3710 4634 3738 4639
rect 3374 4578 3402 4583
rect 3262 4577 3402 4578
rect 3262 4551 3375 4577
rect 3401 4551 3402 4577
rect 3262 4550 3402 4551
rect 3374 4545 3402 4550
rect 3710 4185 3738 4606
rect 3710 4159 3711 4185
rect 3737 4159 3738 4185
rect 3710 4153 3738 4159
rect 3766 4130 3794 5279
rect 3934 5305 3962 5311
rect 3934 5279 3935 5305
rect 3961 5279 3962 5305
rect 3934 5250 3962 5279
rect 3934 5217 3962 5222
rect 4046 5194 4074 5951
rect 4046 5161 4074 5166
rect 4102 5250 4130 5255
rect 4214 5250 4242 6286
rect 4382 6258 4410 6398
rect 4438 6393 4466 6398
rect 4606 6426 4634 6510
rect 4606 6379 4634 6398
rect 4270 6230 4410 6258
rect 4270 6145 4298 6230
rect 4270 6119 4271 6145
rect 4297 6119 4298 6145
rect 4270 6113 4298 6119
rect 4326 6146 4354 6151
rect 4270 5754 4298 5759
rect 4326 5754 4354 6118
rect 4494 6145 4522 6151
rect 4494 6119 4495 6145
rect 4521 6119 4522 6145
rect 4270 5753 4354 5754
rect 4270 5727 4271 5753
rect 4297 5727 4354 5753
rect 4270 5726 4354 5727
rect 4382 6090 4410 6095
rect 4270 5721 4298 5726
rect 4130 5222 4242 5250
rect 4270 5361 4298 5367
rect 4270 5335 4271 5361
rect 4297 5335 4298 5361
rect 4270 5250 4298 5335
rect 4382 5362 4410 6062
rect 4438 5586 4466 5591
rect 4494 5586 4522 6119
rect 4662 6146 4690 6566
rect 4718 6481 4746 6734
rect 5054 6593 5082 6958
rect 5166 6930 5194 7014
rect 5110 6762 5138 6767
rect 5110 6715 5138 6734
rect 5054 6567 5055 6593
rect 5081 6567 5082 6593
rect 5054 6561 5082 6567
rect 5166 6593 5194 6902
rect 5334 6874 5362 7239
rect 5558 7210 5586 7215
rect 5558 7163 5586 7182
rect 5614 7153 5642 7159
rect 5614 7127 5615 7153
rect 5641 7127 5642 7153
rect 5614 7098 5642 7127
rect 5670 7154 5698 7159
rect 5670 7107 5698 7126
rect 5726 7153 5754 7159
rect 5726 7127 5727 7153
rect 5753 7127 5754 7153
rect 5278 6846 5362 6874
rect 5390 7070 5642 7098
rect 5166 6567 5167 6593
rect 5193 6567 5194 6593
rect 5166 6561 5194 6567
rect 5222 6818 5250 6823
rect 4718 6455 4719 6481
rect 4745 6455 4746 6481
rect 4718 6449 4746 6455
rect 4918 6286 5050 6291
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 4918 6253 5050 6258
rect 5166 6258 5194 6263
rect 4830 6202 4858 6207
rect 4830 6155 4858 6174
rect 5054 6202 5082 6207
rect 4550 5977 4578 5983
rect 4550 5951 4551 5977
rect 4577 5951 4578 5977
rect 4550 5698 4578 5951
rect 4550 5665 4578 5670
rect 4606 5698 4634 5703
rect 4662 5698 4690 6118
rect 4998 6090 5026 6095
rect 4606 5697 4690 5698
rect 4606 5671 4607 5697
rect 4633 5671 4690 5697
rect 4606 5670 4690 5671
rect 4718 6089 5026 6090
rect 4718 6063 4999 6089
rect 5025 6063 5026 6089
rect 4718 6062 5026 6063
rect 4606 5665 4634 5670
rect 4438 5585 4578 5586
rect 4438 5559 4439 5585
rect 4465 5559 4578 5585
rect 4438 5558 4578 5559
rect 4438 5553 4466 5558
rect 4438 5362 4466 5367
rect 4382 5334 4438 5362
rect 3840 5110 3972 5115
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3840 5077 3972 5082
rect 4102 5082 4130 5222
rect 4270 5217 4298 5222
rect 4438 5249 4466 5334
rect 4438 5223 4439 5249
rect 4465 5223 4466 5249
rect 4438 5217 4466 5223
rect 4494 5305 4522 5311
rect 4494 5279 4495 5305
rect 4521 5279 4522 5305
rect 4102 5049 4130 5054
rect 4438 4465 4466 4471
rect 4438 4439 4439 4465
rect 4465 4439 4466 4465
rect 3840 4326 3972 4331
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3840 4293 3972 4298
rect 3766 4102 4018 4130
rect 3654 4017 3682 4023
rect 3766 4018 3794 4023
rect 3654 3991 3655 4017
rect 3681 3991 3682 4017
rect 3094 3761 3122 3766
rect 3374 3822 3626 3850
rect 3374 3793 3402 3822
rect 3374 3767 3375 3793
rect 3401 3767 3402 3793
rect 3038 3738 3066 3743
rect 2814 3065 2954 3066
rect 2814 3039 2815 3065
rect 2841 3039 2954 3065
rect 2814 3038 2954 3039
rect 2982 3737 3066 3738
rect 2982 3711 3039 3737
rect 3065 3711 3066 3737
rect 2982 3710 3066 3711
rect 2982 3345 3010 3710
rect 3038 3705 3066 3710
rect 3150 3738 3178 3743
rect 3150 3691 3178 3710
rect 3206 3625 3234 3631
rect 3206 3599 3207 3625
rect 3233 3599 3234 3625
rect 2982 3319 2983 3345
rect 3009 3319 3010 3345
rect 2142 2954 2170 2959
rect 2142 2169 2170 2926
rect 2814 2954 2842 3038
rect 2814 2921 2842 2926
rect 2590 2897 2618 2903
rect 2590 2871 2591 2897
rect 2617 2871 2618 2897
rect 2590 2842 2618 2871
rect 2982 2842 3010 3319
rect 3038 3514 3066 3519
rect 3038 2953 3066 3486
rect 3094 3458 3122 3463
rect 3094 3411 3122 3430
rect 3094 3066 3122 3071
rect 3094 3019 3122 3038
rect 3206 3065 3234 3599
rect 3206 3039 3207 3065
rect 3233 3039 3234 3065
rect 3038 2927 3039 2953
rect 3065 2927 3066 2953
rect 3038 2921 3066 2927
rect 3150 2897 3178 2903
rect 3150 2871 3151 2897
rect 3177 2871 3178 2897
rect 2590 2814 3066 2842
rect 2478 2618 2506 2623
rect 2478 2225 2506 2590
rect 2926 2618 2954 2623
rect 2926 2571 2954 2590
rect 2590 2562 2618 2567
rect 2590 2515 2618 2534
rect 2982 2562 3010 2567
rect 2982 2505 3010 2534
rect 2982 2479 2983 2505
rect 3009 2479 3010 2505
rect 2982 2473 3010 2479
rect 2762 2366 2894 2371
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2762 2333 2894 2338
rect 2478 2199 2479 2225
rect 2505 2199 2506 2225
rect 2478 2193 2506 2199
rect 2142 2143 2143 2169
rect 2169 2143 2170 2169
rect 2142 2137 2170 2143
rect 3038 2170 3066 2814
rect 3094 2674 3122 2679
rect 3150 2674 3178 2871
rect 3206 2898 3234 3039
rect 3206 2786 3234 2870
rect 3318 2954 3346 2959
rect 3374 2954 3402 3767
rect 3542 3737 3570 3743
rect 3542 3711 3543 3737
rect 3569 3711 3570 3737
rect 3542 3570 3570 3711
rect 3598 3626 3626 3822
rect 3654 3738 3682 3991
rect 3654 3705 3682 3710
rect 3710 4017 3794 4018
rect 3710 3991 3767 4017
rect 3793 3991 3794 4017
rect 3710 3990 3794 3991
rect 3710 3681 3738 3990
rect 3766 3985 3794 3990
rect 3878 4018 3906 4023
rect 3878 3971 3906 3990
rect 3990 3850 4018 4102
rect 4438 4018 4466 4439
rect 4494 4074 4522 5279
rect 4550 5306 4578 5558
rect 4550 5273 4578 5278
rect 4494 4041 4522 4046
rect 4550 4970 4578 4975
rect 4550 4185 4578 4942
rect 4718 4410 4746 6062
rect 4998 6057 5026 6062
rect 4942 5978 4970 5983
rect 4942 5753 4970 5950
rect 4942 5727 4943 5753
rect 4969 5727 4970 5753
rect 4942 5721 4970 5727
rect 4886 5698 4914 5703
rect 4886 5651 4914 5670
rect 4998 5698 5026 5703
rect 4998 5651 5026 5670
rect 5054 5586 5082 6174
rect 5166 6090 5194 6230
rect 5222 6201 5250 6790
rect 5278 6594 5306 6846
rect 5334 6761 5362 6767
rect 5334 6735 5335 6761
rect 5361 6735 5362 6761
rect 5334 6650 5362 6735
rect 5334 6617 5362 6622
rect 5278 6561 5306 6566
rect 5334 6538 5362 6543
rect 5334 6491 5362 6510
rect 5278 6481 5306 6487
rect 5278 6455 5279 6481
rect 5305 6455 5306 6481
rect 5278 6426 5306 6455
rect 5278 6393 5306 6398
rect 5334 6370 5362 6375
rect 5390 6370 5418 7070
rect 5726 7042 5754 7127
rect 5614 7014 5754 7042
rect 5334 6369 5418 6370
rect 5334 6343 5335 6369
rect 5361 6343 5418 6369
rect 5334 6342 5418 6343
rect 5502 6538 5530 6543
rect 5334 6337 5362 6342
rect 5222 6175 5223 6201
rect 5249 6175 5250 6201
rect 5222 6169 5250 6175
rect 5278 6314 5306 6319
rect 5278 6090 5306 6286
rect 5390 6202 5418 6207
rect 5110 6089 5194 6090
rect 5110 6063 5167 6089
rect 5193 6063 5194 6089
rect 5110 6062 5194 6063
rect 5110 5698 5138 6062
rect 5166 6057 5194 6062
rect 5222 6062 5306 6090
rect 5334 6089 5362 6095
rect 5334 6063 5335 6089
rect 5361 6063 5362 6089
rect 5166 5810 5194 5815
rect 5166 5763 5194 5782
rect 5110 5665 5138 5670
rect 5166 5697 5194 5703
rect 5166 5671 5167 5697
rect 5193 5671 5194 5697
rect 5166 5586 5194 5671
rect 5054 5558 5138 5586
rect 4918 5502 5050 5507
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 4918 5469 5050 5474
rect 4774 5362 4802 5367
rect 4774 5315 4802 5334
rect 4830 5361 4858 5367
rect 4830 5335 4831 5361
rect 4857 5335 4858 5361
rect 4830 5306 4858 5335
rect 4774 5194 4802 5199
rect 4774 4577 4802 5166
rect 4830 4633 4858 5278
rect 4942 5306 4970 5311
rect 4942 5259 4970 5278
rect 5110 5305 5138 5558
rect 5166 5553 5194 5558
rect 5110 5279 5111 5305
rect 5137 5279 5138 5305
rect 5110 5273 5138 5279
rect 5222 5306 5250 6062
rect 5278 5978 5306 5983
rect 5278 5931 5306 5950
rect 5334 5474 5362 6063
rect 5334 5441 5362 5446
rect 5222 5273 5250 5278
rect 5334 5362 5362 5367
rect 4918 4718 5050 4723
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 4918 4685 5050 4690
rect 4830 4607 4831 4633
rect 4857 4607 4858 4633
rect 4830 4601 4858 4607
rect 4774 4551 4775 4577
rect 4801 4551 4802 4577
rect 4774 4545 4802 4551
rect 5334 4521 5362 5334
rect 5390 5250 5418 6174
rect 5502 6090 5530 6510
rect 5558 6425 5586 6431
rect 5558 6399 5559 6425
rect 5585 6399 5586 6425
rect 5558 6314 5586 6399
rect 5558 6281 5586 6286
rect 5558 6090 5586 6095
rect 5502 6089 5586 6090
rect 5502 6063 5559 6089
rect 5585 6063 5586 6089
rect 5502 6062 5586 6063
rect 5558 6057 5586 6062
rect 5614 5698 5642 7014
rect 5782 6986 5810 7630
rect 6230 7602 6258 7607
rect 6174 7574 6230 7602
rect 5996 7462 6128 7467
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 5996 7429 6128 7434
rect 5950 7377 5978 7383
rect 5950 7351 5951 7377
rect 5977 7351 5978 7377
rect 5894 7266 5922 7271
rect 5894 7219 5922 7238
rect 5726 6958 5810 6986
rect 5838 7154 5866 7159
rect 5838 6986 5866 7126
rect 5950 6986 5978 7351
rect 6174 7266 6202 7574
rect 6230 7569 6258 7574
rect 6062 7238 6202 7266
rect 6398 7321 6426 7910
rect 7074 7854 7206 7859
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7074 7821 7206 7826
rect 7910 7769 7938 9198
rect 8582 8386 8610 8391
rect 8152 8246 8284 8251
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8152 8213 8284 8218
rect 8582 8106 8610 8358
rect 8190 8050 8218 8055
rect 8190 8003 8218 8022
rect 8582 8049 8610 8078
rect 8862 8106 8890 8111
rect 8862 8059 8890 8078
rect 8582 8023 8583 8049
rect 8609 8023 8610 8049
rect 8582 8017 8610 8023
rect 8806 8050 8834 8055
rect 7910 7743 7911 7769
rect 7937 7743 7938 7769
rect 7910 7737 7938 7743
rect 8470 7937 8498 7943
rect 8470 7911 8471 7937
rect 8497 7911 8498 7937
rect 6902 7658 6930 7663
rect 6902 7611 6930 7630
rect 7574 7658 7602 7663
rect 6510 7602 6538 7607
rect 6510 7555 6538 7574
rect 6398 7295 6399 7321
rect 6425 7295 6426 7321
rect 6398 7266 6426 7295
rect 6006 7154 6034 7173
rect 6006 7121 6034 7126
rect 5670 6481 5698 6487
rect 5670 6455 5671 6481
rect 5697 6455 5698 6481
rect 5670 6370 5698 6455
rect 5726 6370 5754 6958
rect 5838 6953 5866 6958
rect 5894 6958 5978 6986
rect 6062 6985 6090 7238
rect 6398 7233 6426 7238
rect 7238 7266 7266 7271
rect 7238 7219 7266 7238
rect 7294 7265 7322 7271
rect 7294 7239 7295 7265
rect 7321 7239 7322 7265
rect 6230 7209 6258 7215
rect 6230 7183 6231 7209
rect 6257 7183 6258 7209
rect 6062 6959 6063 6985
rect 6089 6959 6090 6985
rect 5838 6873 5866 6879
rect 5838 6847 5839 6873
rect 5865 6847 5866 6873
rect 5782 6706 5810 6711
rect 5782 6593 5810 6678
rect 5782 6567 5783 6593
rect 5809 6567 5810 6593
rect 5782 6561 5810 6567
rect 5782 6370 5810 6375
rect 5726 6369 5810 6370
rect 5726 6343 5783 6369
rect 5809 6343 5810 6369
rect 5726 6342 5810 6343
rect 5670 6337 5698 6342
rect 5782 6337 5810 6342
rect 5838 6258 5866 6847
rect 5894 6481 5922 6958
rect 6062 6953 6090 6959
rect 6118 7153 6146 7159
rect 6118 7127 6119 7153
rect 6145 7127 6146 7153
rect 5950 6874 5978 6879
rect 5950 6827 5978 6846
rect 6062 6762 6090 6781
rect 6118 6762 6146 7127
rect 6174 6874 6202 6879
rect 6174 6827 6202 6846
rect 6118 6734 6202 6762
rect 6062 6729 6090 6734
rect 5996 6678 6128 6683
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 5996 6645 6128 6650
rect 6174 6594 6202 6734
rect 6174 6561 6202 6566
rect 6230 6538 6258 7183
rect 6454 7210 6482 7215
rect 6454 7042 6482 7182
rect 7014 7209 7042 7215
rect 7014 7183 7015 7209
rect 7041 7183 7042 7209
rect 6286 7014 6482 7042
rect 6678 7154 6706 7159
rect 6286 6873 6314 7014
rect 6678 6986 6706 7126
rect 6902 6986 6930 6991
rect 6454 6985 6930 6986
rect 6454 6959 6679 6985
rect 6705 6959 6903 6985
rect 6929 6959 6930 6985
rect 6454 6958 6930 6959
rect 6286 6847 6287 6873
rect 6313 6847 6314 6873
rect 6286 6841 6314 6847
rect 6398 6873 6426 6879
rect 6398 6847 6399 6873
rect 6425 6847 6426 6873
rect 6398 6538 6426 6847
rect 6230 6510 6426 6538
rect 5894 6455 5895 6481
rect 5921 6455 5922 6481
rect 5894 6449 5922 6455
rect 6006 6482 6034 6487
rect 5838 6225 5866 6230
rect 5726 6146 5754 6151
rect 5950 6146 5978 6151
rect 5726 6145 5978 6146
rect 5726 6119 5727 6145
rect 5753 6119 5951 6145
rect 5977 6119 5978 6145
rect 5726 6118 5978 6119
rect 5726 6113 5754 6118
rect 5950 6090 5978 6118
rect 5950 6057 5978 6062
rect 5726 6034 5754 6039
rect 5726 5810 5754 6006
rect 5894 5978 5922 5983
rect 5894 5931 5922 5950
rect 6006 5978 6034 6454
rect 6174 6426 6202 6431
rect 6174 6379 6202 6398
rect 6006 5945 6034 5950
rect 6062 6314 6090 6319
rect 6286 6314 6314 6510
rect 6454 6482 6482 6958
rect 6678 6953 6706 6958
rect 6902 6953 6930 6958
rect 6510 6874 6538 6879
rect 6510 6817 6538 6846
rect 6510 6791 6511 6817
rect 6537 6791 6538 6817
rect 6510 6785 6538 6791
rect 6566 6873 6594 6879
rect 6566 6847 6567 6873
rect 6593 6847 6594 6873
rect 6342 6454 6482 6482
rect 6566 6594 6594 6847
rect 6958 6874 6986 6879
rect 7014 6874 7042 7183
rect 7126 7210 7154 7215
rect 7126 7163 7154 7182
rect 7074 7070 7206 7075
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7074 7037 7206 7042
rect 6958 6873 7098 6874
rect 6958 6847 6959 6873
rect 6985 6847 7098 6873
rect 6958 6846 7098 6847
rect 6958 6841 6986 6846
rect 6342 6425 6370 6454
rect 6342 6399 6343 6425
rect 6369 6399 6370 6425
rect 6342 6370 6370 6399
rect 6342 6342 6426 6370
rect 6286 6286 6370 6314
rect 6062 6034 6090 6286
rect 6062 5978 6090 6006
rect 6286 6033 6314 6039
rect 6286 6007 6287 6033
rect 6313 6007 6314 6033
rect 6230 5978 6258 5983
rect 6062 5977 6258 5978
rect 6062 5951 6063 5977
rect 6089 5951 6231 5977
rect 6257 5951 6258 5977
rect 6062 5950 6258 5951
rect 6062 5945 6090 5950
rect 6230 5945 6258 5950
rect 5996 5894 6128 5899
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 5996 5861 6128 5866
rect 6286 5810 6314 6007
rect 5726 5809 5922 5810
rect 5726 5783 5727 5809
rect 5753 5783 5922 5809
rect 5726 5782 5922 5783
rect 5726 5777 5754 5782
rect 5558 5670 5642 5698
rect 5446 5250 5474 5255
rect 5390 5222 5446 5250
rect 5334 4495 5335 4521
rect 5361 4495 5362 4521
rect 4830 4410 4858 4415
rect 4718 4409 4858 4410
rect 4718 4383 4831 4409
rect 4857 4383 4858 4409
rect 4718 4382 4858 4383
rect 4830 4377 4858 4382
rect 4550 4159 4551 4185
rect 4577 4159 4578 4185
rect 4438 3985 4466 3990
rect 3990 3849 4074 3850
rect 3990 3823 3991 3849
rect 4017 3823 4074 3849
rect 3990 3822 4074 3823
rect 3990 3817 4018 3822
rect 3710 3655 3711 3681
rect 3737 3655 3738 3681
rect 3710 3626 3738 3655
rect 3822 3738 3850 3743
rect 3822 3626 3850 3710
rect 3598 3598 3738 3626
rect 3766 3625 3850 3626
rect 3766 3599 3823 3625
rect 3849 3599 3850 3625
rect 3766 3598 3850 3599
rect 3542 3542 3682 3570
rect 3318 2953 3402 2954
rect 3318 2927 3319 2953
rect 3345 2927 3402 2953
rect 3318 2926 3402 2927
rect 3430 3345 3458 3351
rect 3430 3319 3431 3345
rect 3457 3319 3458 3345
rect 3206 2758 3290 2786
rect 3094 2673 3178 2674
rect 3094 2647 3095 2673
rect 3121 2647 3178 2673
rect 3094 2646 3178 2647
rect 3094 2641 3122 2646
rect 3262 2505 3290 2758
rect 3318 2674 3346 2926
rect 3318 2641 3346 2646
rect 3430 2562 3458 3319
rect 3654 3346 3682 3542
rect 3766 3458 3794 3598
rect 3822 3593 3850 3598
rect 3840 3542 3972 3547
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3840 3509 3972 3514
rect 3766 3430 3906 3458
rect 3654 3299 3682 3318
rect 3486 3066 3514 3071
rect 3486 3019 3514 3038
rect 3710 2954 3738 2959
rect 3430 2561 3570 2562
rect 3430 2535 3431 2561
rect 3457 2535 3570 2561
rect 3430 2534 3570 2535
rect 3430 2529 3458 2534
rect 3262 2479 3263 2505
rect 3289 2479 3290 2505
rect 3262 2473 3290 2479
rect 3094 2170 3122 2175
rect 3038 2142 3094 2170
rect 3094 2137 3122 2142
rect 3542 2113 3570 2534
rect 3542 2087 3543 2113
rect 3569 2087 3570 2113
rect 3542 2081 3570 2087
rect 3710 1833 3738 2926
rect 3822 2953 3850 2959
rect 3822 2927 3823 2953
rect 3849 2927 3850 2953
rect 3766 2898 3794 2903
rect 3822 2898 3850 2927
rect 3794 2870 3850 2898
rect 3878 2897 3906 3430
rect 3878 2871 3879 2897
rect 3905 2871 3906 2897
rect 3766 2170 3794 2870
rect 3878 2865 3906 2871
rect 3934 3346 3962 3351
rect 3934 2953 3962 3318
rect 4046 3345 4074 3822
rect 4046 3319 4047 3345
rect 4073 3319 4074 3345
rect 4046 3313 4074 3319
rect 4270 3401 4298 3407
rect 4270 3375 4271 3401
rect 4297 3375 4298 3401
rect 4158 3289 4186 3295
rect 4158 3263 4159 3289
rect 4185 3263 4186 3289
rect 4158 3066 4186 3263
rect 4214 3290 4242 3295
rect 4214 3233 4242 3262
rect 4214 3207 4215 3233
rect 4241 3207 4242 3233
rect 4214 3201 4242 3207
rect 4270 3122 4298 3375
rect 4270 3089 4298 3094
rect 4382 3345 4410 3351
rect 4550 3346 4578 4159
rect 5222 4129 5250 4135
rect 5222 4103 5223 4129
rect 5249 4103 5250 4129
rect 4942 4074 4970 4079
rect 4942 4027 4970 4046
rect 5222 4018 5250 4103
rect 5334 4130 5362 4495
rect 5390 4466 5418 4471
rect 5390 4419 5418 4438
rect 5390 4130 5418 4135
rect 5334 4129 5418 4130
rect 5334 4103 5391 4129
rect 5417 4103 5418 4129
rect 5334 4102 5418 4103
rect 5222 3985 5250 3990
rect 4918 3934 5050 3939
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 4918 3901 5050 3906
rect 5390 3626 5418 4102
rect 5446 3793 5474 5222
rect 5558 4578 5586 5670
rect 5894 5641 5922 5782
rect 6286 5777 6314 5782
rect 5894 5615 5895 5641
rect 5921 5615 5922 5641
rect 5894 5609 5922 5615
rect 5950 5698 5978 5703
rect 5614 5585 5642 5591
rect 5614 5559 5615 5585
rect 5641 5559 5642 5585
rect 5614 5362 5642 5559
rect 5670 5586 5698 5591
rect 5670 5539 5698 5558
rect 5950 5530 5978 5670
rect 6062 5698 6090 5703
rect 6342 5698 6370 6286
rect 6398 6089 6426 6342
rect 6398 6063 6399 6089
rect 6425 6063 6426 6089
rect 6398 6057 6426 6063
rect 6566 6090 6594 6566
rect 6902 6761 6930 6767
rect 6902 6735 6903 6761
rect 6929 6735 6930 6761
rect 6790 6146 6818 6151
rect 6902 6146 6930 6735
rect 6958 6650 6986 6655
rect 6958 6370 6986 6622
rect 7070 6538 7098 6846
rect 7294 6650 7322 7239
rect 7574 7266 7602 7630
rect 8414 7658 8442 7663
rect 8414 7611 8442 7630
rect 8152 7462 8284 7467
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8152 7429 8284 7434
rect 7574 7265 7658 7266
rect 7574 7239 7575 7265
rect 7601 7239 7658 7265
rect 7574 7238 7658 7239
rect 7574 7233 7602 7238
rect 7518 7210 7546 7215
rect 7294 6617 7322 6622
rect 7406 7153 7434 7159
rect 7406 7127 7407 7153
rect 7433 7127 7434 7153
rect 7406 6538 7434 7127
rect 7070 6510 7378 6538
rect 6958 6337 6986 6342
rect 7014 6482 7042 6487
rect 6790 6145 6874 6146
rect 6790 6119 6791 6145
rect 6817 6119 6874 6145
rect 6790 6118 6874 6119
rect 6790 6113 6818 6118
rect 6566 6057 6594 6062
rect 6062 5697 6370 5698
rect 6062 5671 6063 5697
rect 6089 5671 6343 5697
rect 6369 5671 6370 5697
rect 6062 5670 6370 5671
rect 6062 5665 6090 5670
rect 5614 5329 5642 5334
rect 5894 5502 5950 5530
rect 5726 5026 5754 5031
rect 5726 4913 5754 4998
rect 5726 4887 5727 4913
rect 5753 4887 5754 4913
rect 5614 4578 5642 4583
rect 5558 4577 5642 4578
rect 5558 4551 5615 4577
rect 5641 4551 5642 4577
rect 5558 4550 5642 4551
rect 5614 4545 5642 4550
rect 5726 4522 5754 4887
rect 5894 4914 5922 5502
rect 5950 5497 5978 5502
rect 6174 5586 6202 5591
rect 6174 5362 6202 5558
rect 6230 5585 6258 5591
rect 6230 5559 6231 5585
rect 6257 5559 6258 5585
rect 6230 5530 6258 5559
rect 6230 5497 6258 5502
rect 6174 5334 6258 5362
rect 6174 5249 6202 5255
rect 6174 5223 6175 5249
rect 6201 5223 6202 5249
rect 5996 5110 6128 5115
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 5996 5077 6128 5082
rect 6174 5026 6202 5223
rect 6174 4993 6202 4998
rect 6230 5025 6258 5334
rect 6230 4999 6231 5025
rect 6257 4999 6258 5025
rect 6230 4993 6258 4999
rect 6118 4970 6146 4975
rect 5950 4914 5978 4919
rect 5894 4913 5978 4914
rect 5894 4887 5951 4913
rect 5977 4887 5978 4913
rect 5894 4886 5978 4887
rect 6118 4914 6146 4942
rect 6118 4886 6202 4914
rect 5950 4881 5978 4886
rect 6062 4857 6090 4863
rect 6062 4831 6063 4857
rect 6089 4831 6090 4857
rect 5782 4522 5810 4527
rect 5726 4521 5810 4522
rect 5726 4495 5783 4521
rect 5809 4495 5810 4521
rect 5726 4494 5810 4495
rect 5782 4489 5810 4494
rect 5894 4466 5922 4471
rect 5894 4410 5922 4438
rect 6062 4410 6090 4831
rect 5894 4382 6090 4410
rect 5894 4242 5922 4382
rect 5996 4326 6128 4331
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 5996 4293 6128 4298
rect 5950 4242 5978 4247
rect 5894 4241 5978 4242
rect 5894 4215 5951 4241
rect 5977 4215 5978 4241
rect 5894 4214 5978 4215
rect 5950 4209 5978 4214
rect 6006 4130 6034 4135
rect 5446 3767 5447 3793
rect 5473 3767 5474 3793
rect 5446 3761 5474 3767
rect 5502 4074 5530 4079
rect 5502 3737 5530 4046
rect 5894 4073 5922 4079
rect 5894 4047 5895 4073
rect 5921 4047 5922 4073
rect 5894 4018 5922 4047
rect 5894 3985 5922 3990
rect 5502 3711 5503 3737
rect 5529 3711 5530 3737
rect 5502 3705 5530 3711
rect 6006 3681 6034 4102
rect 6174 3737 6202 4886
rect 6286 4690 6314 5670
rect 6342 5665 6370 5670
rect 6846 5697 6874 6118
rect 6902 6113 6930 6118
rect 6958 6146 6986 6151
rect 7014 6146 7042 6454
rect 7294 6426 7322 6431
rect 7238 6398 7294 6426
rect 7126 6370 7154 6389
rect 7126 6337 7154 6342
rect 7074 6286 7206 6291
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7074 6253 7206 6258
rect 6958 6145 7042 6146
rect 6958 6119 6959 6145
rect 6985 6119 7042 6145
rect 6958 6118 7042 6119
rect 6958 6113 6986 6118
rect 6846 5671 6847 5697
rect 6873 5671 6874 5697
rect 6734 5642 6762 5647
rect 6734 5595 6762 5614
rect 6342 5586 6370 5591
rect 6342 4913 6370 5558
rect 6342 4887 6343 4913
rect 6369 4887 6370 4913
rect 6342 4881 6370 4887
rect 6734 5418 6762 5423
rect 6342 4802 6370 4807
rect 6734 4802 6762 5390
rect 6846 4914 6874 5671
rect 7182 5866 7210 5871
rect 7182 5697 7210 5838
rect 7182 5671 7183 5697
rect 7209 5671 7210 5697
rect 7182 5665 7210 5671
rect 7070 5642 7098 5647
rect 7070 5595 7098 5614
rect 7074 5502 7206 5507
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7074 5469 7206 5474
rect 7182 5418 7210 5423
rect 7182 4970 7210 5390
rect 7238 5306 7266 6398
rect 7294 6379 7322 6398
rect 7350 6370 7378 6510
rect 7406 6505 7434 6510
rect 7462 6370 7490 6375
rect 7350 6369 7490 6370
rect 7350 6343 7463 6369
rect 7489 6343 7490 6369
rect 7350 6342 7490 6343
rect 7350 6258 7378 6263
rect 7294 5754 7322 5759
rect 7294 5707 7322 5726
rect 7350 5697 7378 6230
rect 7350 5671 7351 5697
rect 7377 5671 7378 5697
rect 7350 5665 7378 5671
rect 7406 5642 7434 6342
rect 7462 6337 7490 6342
rect 7406 5609 7434 5614
rect 7462 5586 7490 5591
rect 7518 5586 7546 7182
rect 7462 5585 7546 5586
rect 7462 5559 7463 5585
rect 7489 5559 7546 5585
rect 7462 5558 7546 5559
rect 7630 6481 7658 7238
rect 7966 7210 7994 7215
rect 7966 7163 7994 7182
rect 8414 6874 8442 6879
rect 8414 6827 8442 6846
rect 7910 6762 7938 6767
rect 7910 6715 7938 6734
rect 8152 6678 8284 6683
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8152 6645 8284 6650
rect 8022 6538 8050 6543
rect 8022 6491 8050 6510
rect 7630 6455 7631 6481
rect 7657 6455 7658 6481
rect 7630 5697 7658 6455
rect 8470 6482 8498 7911
rect 8806 7770 8834 8022
rect 9230 7854 9362 7859
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9230 7821 9362 7826
rect 8806 7769 9058 7770
rect 8806 7743 8807 7769
rect 8833 7743 9058 7769
rect 8806 7742 9058 7743
rect 8806 7737 8834 7742
rect 8806 7601 8834 7607
rect 8806 7575 8807 7601
rect 8833 7575 8834 7601
rect 8470 6449 8498 6454
rect 8694 7545 8722 7551
rect 8694 7519 8695 7545
rect 8721 7519 8722 7545
rect 8694 6761 8722 7519
rect 8750 7266 8778 7271
rect 8750 6985 8778 7238
rect 8750 6959 8751 6985
rect 8777 6959 8778 6985
rect 8750 6953 8778 6959
rect 8694 6735 8695 6761
rect 8721 6735 8722 6761
rect 8694 6426 8722 6735
rect 8694 6393 8722 6398
rect 8638 6146 8666 6151
rect 7966 6090 7994 6095
rect 7630 5671 7631 5697
rect 7657 5671 7658 5697
rect 7462 5553 7490 5558
rect 7462 5306 7490 5311
rect 7238 5278 7462 5306
rect 7182 4942 7322 4970
rect 7126 4914 7154 4919
rect 6846 4913 7266 4914
rect 6846 4887 6847 4913
rect 6873 4887 7127 4913
rect 7153 4887 7266 4913
rect 6846 4886 7266 4887
rect 6846 4881 6874 4886
rect 7126 4881 7154 4886
rect 6958 4802 6986 4807
rect 6342 4801 6594 4802
rect 6342 4775 6343 4801
rect 6369 4775 6594 4801
rect 6342 4774 6594 4775
rect 6734 4801 6986 4802
rect 6734 4775 6959 4801
rect 6985 4775 6986 4801
rect 6734 4774 6986 4775
rect 6342 4769 6370 4774
rect 6286 4662 6482 4690
rect 6286 4130 6314 4135
rect 6286 4073 6314 4102
rect 6286 4047 6287 4073
rect 6313 4047 6314 4073
rect 6286 4041 6314 4047
rect 6398 4073 6426 4079
rect 6398 4047 6399 4073
rect 6425 4047 6426 4073
rect 6174 3711 6175 3737
rect 6201 3711 6202 3737
rect 6174 3705 6202 3711
rect 6342 4017 6370 4023
rect 6342 3991 6343 4017
rect 6369 3991 6370 4017
rect 6006 3655 6007 3681
rect 6033 3655 6034 3681
rect 6006 3649 6034 3655
rect 5390 3598 5530 3626
rect 5278 3402 5306 3407
rect 4606 3346 4634 3351
rect 4382 3319 4383 3345
rect 4409 3319 4410 3345
rect 4158 3033 4186 3038
rect 4382 3010 4410 3319
rect 4438 3345 4634 3346
rect 4438 3319 4607 3345
rect 4633 3319 4634 3345
rect 4438 3318 4634 3319
rect 4438 3065 4466 3318
rect 4606 3313 4634 3318
rect 4998 3290 5026 3295
rect 4998 3243 5026 3262
rect 4918 3150 5050 3155
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 4918 3117 5050 3122
rect 4438 3039 4439 3065
rect 4465 3039 4466 3065
rect 4438 3033 4466 3039
rect 5222 3066 5250 3071
rect 5222 3019 5250 3038
rect 4382 2977 4410 2982
rect 4998 3010 5026 3015
rect 4998 2963 5026 2982
rect 5278 3009 5306 3374
rect 5278 2983 5279 3009
rect 5305 2983 5306 3009
rect 5278 2977 5306 2983
rect 3934 2927 3935 2953
rect 3961 2927 3962 2953
rect 3934 2898 3962 2927
rect 3990 2898 4018 2903
rect 3934 2870 3990 2898
rect 3990 2865 4018 2870
rect 4998 2897 5026 2903
rect 4998 2871 4999 2897
rect 5025 2871 5026 2897
rect 4046 2842 4074 2847
rect 3840 2758 3972 2763
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3840 2725 3972 2730
rect 3878 2674 3906 2679
rect 3822 2170 3850 2175
rect 3766 2169 3850 2170
rect 3766 2143 3823 2169
rect 3849 2143 3850 2169
rect 3766 2142 3850 2143
rect 3822 2137 3850 2142
rect 3766 2058 3794 2063
rect 3878 2058 3906 2646
rect 3990 2226 4018 2231
rect 4046 2226 4074 2814
rect 4886 2842 4914 2847
rect 4886 2795 4914 2814
rect 4942 2617 4970 2623
rect 4942 2591 4943 2617
rect 4969 2591 4970 2617
rect 3990 2225 4074 2226
rect 3990 2199 3991 2225
rect 4017 2199 4074 2225
rect 3990 2198 4074 2199
rect 4102 2561 4130 2567
rect 4102 2535 4103 2561
rect 4129 2535 4130 2561
rect 3990 2193 4018 2198
rect 3934 2170 3962 2175
rect 3934 2123 3962 2142
rect 3766 2057 3906 2058
rect 3766 2031 3767 2057
rect 3793 2031 3906 2057
rect 3766 2030 3906 2031
rect 3766 2025 3794 2030
rect 3840 1974 3972 1979
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3840 1941 3972 1946
rect 3710 1807 3711 1833
rect 3737 1807 3738 1833
rect 3710 1801 3738 1807
rect 1918 1751 1919 1777
rect 1945 1751 1946 1777
rect 1918 1745 1946 1751
rect 4102 1778 4130 2535
rect 4326 2562 4354 2567
rect 4326 2515 4354 2534
rect 4774 2561 4802 2567
rect 4774 2535 4775 2561
rect 4801 2535 4802 2561
rect 4718 2450 4746 2455
rect 4718 2403 4746 2422
rect 4774 2282 4802 2535
rect 4942 2450 4970 2591
rect 4998 2618 5026 2871
rect 5502 2897 5530 3598
rect 5996 3542 6128 3547
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 5996 3509 6128 3514
rect 6286 3458 6314 3463
rect 6342 3458 6370 3991
rect 6286 3457 6370 3458
rect 6286 3431 6287 3457
rect 6313 3431 6370 3457
rect 6286 3430 6370 3431
rect 6286 3425 6314 3430
rect 6062 3402 6090 3407
rect 6062 3355 6090 3374
rect 6398 3346 6426 4047
rect 6454 3457 6482 4662
rect 6454 3431 6455 3457
rect 6481 3431 6482 3457
rect 6454 3425 6482 3431
rect 6398 3318 6482 3346
rect 6398 3233 6426 3239
rect 6398 3207 6399 3233
rect 6425 3207 6426 3233
rect 6398 3066 6426 3207
rect 6342 3038 6426 3066
rect 5502 2871 5503 2897
rect 5529 2871 5530 2897
rect 5502 2865 5530 2871
rect 6230 2898 6258 2903
rect 5996 2758 6128 2763
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 5996 2725 6128 2730
rect 4998 2585 5026 2590
rect 6006 2618 6034 2623
rect 6006 2571 6034 2590
rect 4942 2422 5250 2450
rect 4918 2366 5050 2371
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 4918 2333 5050 2338
rect 5110 2338 5138 2343
rect 4774 2249 4802 2254
rect 5110 2281 5138 2310
rect 5110 2255 5111 2281
rect 5137 2255 5138 2281
rect 5110 2249 5138 2255
rect 5222 2282 5250 2422
rect 5614 2282 5642 2287
rect 5222 2281 5474 2282
rect 5222 2255 5223 2281
rect 5249 2255 5474 2281
rect 5222 2254 5474 2255
rect 5222 2249 5250 2254
rect 5446 2225 5474 2254
rect 5446 2199 5447 2225
rect 5473 2199 5474 2225
rect 5446 2193 5474 2199
rect 5614 2225 5642 2254
rect 6230 2281 6258 2870
rect 6230 2255 6231 2281
rect 6257 2255 6258 2281
rect 6230 2249 6258 2255
rect 6342 2282 6370 3038
rect 6398 2954 6426 2959
rect 6398 2561 6426 2926
rect 6398 2535 6399 2561
rect 6425 2535 6426 2561
rect 6398 2529 6426 2535
rect 6454 2450 6482 3318
rect 6566 3009 6594 4774
rect 6958 4466 6986 4774
rect 7074 4718 7206 4723
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7074 4685 7206 4690
rect 6958 4433 6986 4438
rect 6734 4186 6930 4214
rect 6734 4185 6762 4186
rect 6734 4159 6735 4185
rect 6761 4159 6762 4185
rect 6734 4130 6762 4159
rect 6846 4130 6874 4135
rect 6734 4097 6762 4102
rect 6790 4129 6874 4130
rect 6790 4103 6847 4129
rect 6873 4103 6874 4129
rect 6790 4102 6874 4103
rect 6566 2983 6567 3009
rect 6593 2983 6594 3009
rect 6566 2977 6594 2983
rect 6790 3401 6818 4102
rect 6846 4097 6874 4102
rect 6790 3375 6791 3401
rect 6817 3375 6818 3401
rect 6454 2417 6482 2422
rect 6678 2562 6706 2567
rect 5614 2199 5615 2225
rect 5641 2199 5642 2225
rect 5614 2193 5642 2199
rect 5278 2170 5306 2175
rect 5278 2123 5306 2142
rect 6342 2169 6370 2254
rect 6342 2143 6343 2169
rect 6369 2143 6370 2169
rect 6342 2137 6370 2143
rect 6622 2282 6650 2287
rect 6622 2170 6650 2254
rect 5996 1974 6128 1979
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 5996 1941 6128 1946
rect 6622 1889 6650 2142
rect 6622 1863 6623 1889
rect 6649 1863 6650 1889
rect 6622 1857 6650 1863
rect 6678 2114 6706 2534
rect 6734 2338 6762 2343
rect 6790 2338 6818 3375
rect 6902 3345 6930 4186
rect 7238 4129 7266 4886
rect 7294 4857 7322 4942
rect 7294 4831 7295 4857
rect 7321 4831 7322 4857
rect 7294 4214 7322 4831
rect 7294 4186 7434 4214
rect 7238 4103 7239 4129
rect 7265 4103 7266 4129
rect 7238 4097 7266 4103
rect 7014 4017 7042 4023
rect 7014 3991 7015 4017
rect 7041 3991 7042 4017
rect 6902 3319 6903 3345
rect 6929 3319 6930 3345
rect 6902 3234 6930 3319
rect 6846 3206 6930 3234
rect 6958 3737 6986 3743
rect 6958 3711 6959 3737
rect 6985 3711 6986 3737
rect 6958 3402 6986 3711
rect 6846 2562 6874 3206
rect 6958 3122 6986 3374
rect 6846 2529 6874 2534
rect 6902 3094 6986 3122
rect 7014 3514 7042 3991
rect 7350 4017 7378 4023
rect 7350 3991 7351 4017
rect 7377 3991 7378 4017
rect 7074 3934 7206 3939
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7074 3901 7206 3906
rect 7350 3850 7378 3991
rect 7350 3817 7378 3822
rect 7406 3849 7434 4186
rect 7406 3823 7407 3849
rect 7433 3823 7434 3849
rect 6902 2561 6930 3094
rect 6958 2954 6986 2959
rect 6958 2907 6986 2926
rect 6958 2786 6986 2791
rect 6958 2617 6986 2758
rect 6958 2591 6959 2617
rect 6985 2591 6986 2617
rect 6958 2585 6986 2591
rect 6902 2535 6903 2561
rect 6929 2535 6930 2561
rect 6902 2529 6930 2535
rect 7014 2561 7042 3486
rect 7070 3794 7098 3799
rect 7070 3457 7098 3766
rect 7294 3626 7322 3631
rect 7070 3431 7071 3457
rect 7097 3431 7098 3457
rect 7070 3425 7098 3431
rect 7238 3625 7322 3626
rect 7238 3599 7295 3625
rect 7321 3599 7322 3625
rect 7238 3598 7322 3599
rect 7074 3150 7206 3155
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7074 3117 7206 3122
rect 7238 2786 7266 3598
rect 7294 3593 7322 3598
rect 7294 3514 7322 3519
rect 7322 3486 7378 3514
rect 7294 3481 7322 3486
rect 7350 3345 7378 3486
rect 7350 3319 7351 3345
rect 7377 3319 7378 3345
rect 7350 3313 7378 3319
rect 7406 3010 7434 3823
rect 7462 3794 7490 5278
rect 7574 4914 7602 4919
rect 7630 4914 7658 5671
rect 7910 5977 7938 5983
rect 7910 5951 7911 5977
rect 7937 5951 7938 5977
rect 7854 5642 7882 5647
rect 7854 5361 7882 5614
rect 7910 5586 7938 5951
rect 7910 5553 7938 5558
rect 7910 5418 7938 5423
rect 7966 5418 7994 6062
rect 8358 6089 8386 6095
rect 8358 6063 8359 6089
rect 8385 6063 8386 6089
rect 8022 6034 8050 6039
rect 8022 5753 8050 6006
rect 8152 5894 8284 5899
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8152 5861 8284 5866
rect 8358 5810 8386 6063
rect 8638 6089 8666 6118
rect 8638 6063 8639 6089
rect 8665 6063 8666 6089
rect 8638 6057 8666 6063
rect 8750 6034 8778 6039
rect 8750 5987 8778 6006
rect 8358 5777 8386 5782
rect 8750 5810 8778 5815
rect 8022 5727 8023 5753
rect 8049 5727 8050 5753
rect 8022 5721 8050 5727
rect 7910 5417 7994 5418
rect 7910 5391 7911 5417
rect 7937 5391 7994 5417
rect 7910 5390 7994 5391
rect 8750 5417 8778 5782
rect 8806 5754 8834 7575
rect 9030 7321 9058 7742
rect 9086 7658 9114 7663
rect 9114 7630 9170 7658
rect 9086 7625 9114 7630
rect 9030 7295 9031 7321
rect 9057 7295 9058 7321
rect 9030 7289 9058 7295
rect 8862 6874 8890 6893
rect 8890 6846 8946 6874
rect 8862 6841 8890 6846
rect 8918 6538 8946 6846
rect 9086 6538 9114 6543
rect 8918 6537 9114 6538
rect 8918 6511 9087 6537
rect 9113 6511 9114 6537
rect 8918 6510 9114 6511
rect 9086 6505 9114 6510
rect 8806 5721 8834 5726
rect 8862 6089 8890 6095
rect 8862 6063 8863 6089
rect 8889 6063 8890 6089
rect 8750 5391 8751 5417
rect 8777 5391 8778 5417
rect 7910 5385 7938 5390
rect 8750 5385 8778 5391
rect 8862 5417 8890 6063
rect 8862 5391 8863 5417
rect 8889 5391 8890 5417
rect 8862 5385 8890 5391
rect 8918 6089 8946 6095
rect 8918 6063 8919 6089
rect 8945 6063 8946 6089
rect 7854 5335 7855 5361
rect 7881 5335 7882 5361
rect 7854 5329 7882 5335
rect 8190 5362 8218 5367
rect 8190 5315 8218 5334
rect 8134 5306 8162 5311
rect 8134 5259 8162 5278
rect 8302 5306 8330 5311
rect 8694 5306 8722 5311
rect 8302 5305 8386 5306
rect 8302 5279 8303 5305
rect 8329 5279 8386 5305
rect 8302 5278 8386 5279
rect 8302 5273 8330 5278
rect 7910 5194 7938 5199
rect 7910 5193 7994 5194
rect 7910 5167 7911 5193
rect 7937 5167 7994 5193
rect 7910 5166 7994 5167
rect 7910 5161 7938 5166
rect 7574 4913 7658 4914
rect 7574 4887 7575 4913
rect 7601 4887 7658 4913
rect 7574 4886 7658 4887
rect 7574 4578 7602 4886
rect 7910 4858 7938 4863
rect 7910 4811 7938 4830
rect 7574 4577 7714 4578
rect 7574 4551 7575 4577
rect 7601 4551 7714 4577
rect 7574 4550 7714 4551
rect 7574 4545 7602 4550
rect 7462 3761 7490 3766
rect 7686 4129 7714 4550
rect 7686 4103 7687 4129
rect 7713 4103 7714 4129
rect 7462 3626 7490 3631
rect 7462 3625 7546 3626
rect 7462 3599 7463 3625
rect 7489 3599 7546 3625
rect 7462 3598 7546 3599
rect 7462 3593 7490 3598
rect 7462 3458 7490 3463
rect 7462 3289 7490 3430
rect 7518 3346 7546 3598
rect 7518 3313 7546 3318
rect 7686 3345 7714 4103
rect 7686 3319 7687 3345
rect 7713 3319 7714 3345
rect 7462 3263 7463 3289
rect 7489 3263 7490 3289
rect 7462 3257 7490 3263
rect 7406 2977 7434 2982
rect 7238 2753 7266 2758
rect 7686 2954 7714 3319
rect 7910 4186 7938 4191
rect 7910 3065 7938 4158
rect 7966 3738 7994 5166
rect 8152 5110 8284 5115
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8152 5077 8284 5082
rect 8302 5026 8330 5031
rect 8302 4466 8330 4998
rect 8358 4578 8386 5278
rect 8358 4545 8386 4550
rect 8638 5305 8722 5306
rect 8638 5279 8695 5305
rect 8721 5279 8722 5305
rect 8638 5278 8722 5279
rect 8358 4466 8386 4471
rect 8302 4438 8358 4466
rect 8152 4326 8284 4331
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8152 4293 8284 4298
rect 8022 4074 8050 4079
rect 8022 4073 8162 4074
rect 8022 4047 8023 4073
rect 8049 4047 8162 4073
rect 8022 4046 8162 4047
rect 8022 4041 8050 4046
rect 8134 3849 8162 4046
rect 8134 3823 8135 3849
rect 8161 3823 8162 3849
rect 8134 3817 8162 3823
rect 8358 3793 8386 4438
rect 8358 3767 8359 3793
rect 8385 3767 8386 3793
rect 8358 3761 8386 3767
rect 8638 3794 8666 5278
rect 8694 5273 8722 5278
rect 8918 5082 8946 6063
rect 9086 5810 9114 5815
rect 9086 5753 9114 5782
rect 9086 5727 9087 5753
rect 9113 5727 9114 5753
rect 9086 5721 9114 5727
rect 9142 5586 9170 7630
rect 9230 7070 9362 7075
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9230 7037 9362 7042
rect 9230 6286 9362 6291
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9230 6253 9362 6258
rect 8918 5049 8946 5054
rect 8974 5558 9170 5586
rect 8974 4970 9002 5558
rect 9230 5502 9362 5507
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9230 5469 9362 5474
rect 8806 4969 9002 4970
rect 8806 4943 8975 4969
rect 9001 4943 9002 4969
rect 8806 4942 9002 4943
rect 8750 4858 8778 4863
rect 8750 4633 8778 4830
rect 8750 4607 8751 4633
rect 8777 4607 8778 4633
rect 8750 4601 8778 4607
rect 8694 4578 8722 4583
rect 8694 4531 8722 4550
rect 8750 3850 8778 3855
rect 8806 3850 8834 4942
rect 8974 4937 9002 4942
rect 9030 5249 9058 5255
rect 9030 5223 9031 5249
rect 9057 5223 9058 5249
rect 8974 4578 9002 4583
rect 9030 4578 9058 5223
rect 9230 4718 9362 4723
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9230 4685 9362 4690
rect 8974 4577 9058 4578
rect 8974 4551 8975 4577
rect 9001 4551 9058 4577
rect 8974 4550 9058 4551
rect 8750 3849 8834 3850
rect 8750 3823 8751 3849
rect 8777 3823 8834 3849
rect 8750 3822 8834 3823
rect 8862 4521 8890 4527
rect 8862 4495 8863 4521
rect 8889 4495 8890 4521
rect 8862 3849 8890 4495
rect 8974 4214 9002 4550
rect 8862 3823 8863 3849
rect 8889 3823 8890 3849
rect 8750 3817 8778 3822
rect 8862 3817 8890 3823
rect 8918 4186 9002 4214
rect 9086 4186 9114 4191
rect 8918 3850 8946 4186
rect 8694 3794 8722 3799
rect 8638 3766 8694 3794
rect 8022 3738 8050 3743
rect 7966 3737 8050 3738
rect 7966 3711 8023 3737
rect 8049 3711 8050 3737
rect 7966 3710 8050 3711
rect 8022 3705 8050 3710
rect 8246 3738 8274 3743
rect 8246 3691 8274 3710
rect 8694 3737 8722 3766
rect 8694 3711 8695 3737
rect 8721 3711 8722 3737
rect 8358 3626 8386 3631
rect 8152 3542 8284 3547
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8152 3509 8284 3514
rect 8022 3346 8050 3351
rect 8022 3299 8050 3318
rect 7910 3039 7911 3065
rect 7937 3039 7938 3065
rect 7910 3033 7938 3039
rect 8078 3066 8106 3071
rect 7014 2535 7015 2561
rect 7041 2535 7042 2561
rect 7014 2529 7042 2535
rect 7126 2618 7154 2623
rect 7126 2561 7154 2590
rect 7126 2535 7127 2561
rect 7153 2535 7154 2561
rect 6846 2450 6874 2455
rect 7126 2450 7154 2535
rect 7686 2562 7714 2926
rect 7686 2529 7714 2534
rect 6874 2422 6986 2450
rect 6846 2403 6874 2422
rect 6762 2310 6818 2338
rect 6734 2305 6762 2310
rect 6958 2225 6986 2422
rect 6958 2199 6959 2225
rect 6985 2199 6986 2225
rect 6958 2193 6986 2199
rect 7014 2422 7154 2450
rect 7238 2506 7266 2511
rect 6174 1834 6202 1839
rect 6174 1787 6202 1806
rect 4102 1745 4130 1750
rect 5054 1778 5082 1783
rect 5054 1731 5082 1750
rect 6622 1778 6650 1783
rect 6622 1721 6650 1750
rect 6678 1777 6706 2086
rect 6678 1751 6679 1777
rect 6705 1751 6706 1777
rect 6678 1745 6706 1751
rect 7014 1777 7042 2422
rect 7074 2366 7206 2371
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7074 2333 7206 2338
rect 7238 2169 7266 2478
rect 7238 2143 7239 2169
rect 7265 2143 7266 2169
rect 7238 2137 7266 2143
rect 7350 2449 7378 2455
rect 7350 2423 7351 2449
rect 7377 2423 7378 2449
rect 7014 1751 7015 1777
rect 7041 1751 7042 1777
rect 7014 1745 7042 1751
rect 7350 1778 7378 2423
rect 8078 1889 8106 3038
rect 8358 2953 8386 3598
rect 8358 2927 8359 2953
rect 8385 2927 8386 2953
rect 8358 2921 8386 2927
rect 8638 3458 8666 3463
rect 8694 3458 8722 3711
rect 8666 3430 8722 3458
rect 8638 2953 8666 3430
rect 8638 2927 8639 2953
rect 8665 2927 8666 2953
rect 8638 2921 8666 2927
rect 8862 2953 8890 2959
rect 8862 2927 8863 2953
rect 8889 2927 8890 2953
rect 8750 2897 8778 2903
rect 8750 2871 8751 2897
rect 8777 2871 8778 2897
rect 8152 2758 8284 2763
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8750 2730 8778 2871
rect 8152 2725 8284 2730
rect 8470 2702 8778 2730
rect 8470 2617 8498 2702
rect 8470 2591 8471 2617
rect 8497 2591 8498 2617
rect 8470 2585 8498 2591
rect 8806 2562 8834 2567
rect 8806 2515 8834 2534
rect 8862 2282 8890 2927
rect 8918 2954 8946 3822
rect 9030 4185 9114 4186
rect 9030 4159 9087 4185
rect 9113 4159 9114 4185
rect 9030 4158 9114 4159
rect 8974 3794 9002 3799
rect 8974 3747 9002 3766
rect 9030 3793 9058 4158
rect 9086 4153 9114 4158
rect 9230 3934 9362 3939
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9230 3901 9362 3906
rect 9030 3767 9031 3793
rect 9057 3767 9058 3793
rect 9030 3626 9058 3767
rect 9142 3738 9170 3743
rect 9142 3691 9170 3710
rect 9030 3593 9058 3598
rect 9086 3402 9114 3407
rect 9086 3401 9170 3402
rect 9086 3375 9087 3401
rect 9113 3375 9170 3401
rect 9086 3374 9170 3375
rect 9086 3369 9114 3374
rect 8918 2953 9114 2954
rect 8918 2927 8919 2953
rect 8945 2927 9114 2953
rect 8918 2926 9114 2927
rect 8918 2921 8946 2926
rect 9086 2617 9114 2926
rect 9086 2591 9087 2617
rect 9113 2591 9114 2617
rect 9086 2585 9114 2591
rect 9142 2618 9170 3374
rect 9230 3150 9362 3155
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9230 3117 9362 3122
rect 9142 2585 9170 2590
rect 9230 2366 9362 2371
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9230 2333 9362 2338
rect 8862 2249 8890 2254
rect 8750 2170 8778 2175
rect 8750 2169 8946 2170
rect 8750 2143 8751 2169
rect 8777 2143 8946 2169
rect 8750 2142 8946 2143
rect 8750 2137 8778 2142
rect 8694 2114 8722 2119
rect 8694 2067 8722 2086
rect 8152 1974 8284 1979
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8152 1941 8284 1946
rect 8078 1863 8079 1889
rect 8105 1863 8106 1889
rect 8078 1857 8106 1863
rect 7350 1745 7378 1750
rect 6622 1695 6623 1721
rect 6649 1695 6650 1721
rect 6622 1689 6650 1695
rect 8806 1721 8834 1727
rect 8806 1695 8807 1721
rect 8833 1695 8834 1721
rect 8806 1610 8834 1695
rect 8918 1721 8946 2142
rect 8918 1695 8919 1721
rect 8945 1695 8946 1721
rect 8918 1689 8946 1695
rect 9086 1721 9114 1727
rect 9086 1695 9087 1721
rect 9113 1695 9114 1721
rect 9086 1610 9114 1695
rect 2762 1582 2894 1587
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2762 1549 2894 1554
rect 4918 1582 5050 1587
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 4918 1549 5050 1554
rect 7074 1582 7206 1587
rect 8806 1582 9114 1610
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7074 1549 7206 1554
rect 966 1241 994 1246
rect 9086 602 9114 1582
rect 9230 1582 9362 1587
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9230 1549 9362 1554
rect 9086 569 9114 574
<< via2 >>
rect 854 8638 882 8666
rect 1684 8245 1712 8246
rect 1684 8219 1685 8245
rect 1685 8219 1711 8245
rect 1711 8219 1712 8245
rect 1684 8218 1712 8219
rect 1736 8245 1764 8246
rect 1736 8219 1737 8245
rect 1737 8219 1763 8245
rect 1763 8219 1764 8245
rect 1736 8218 1764 8219
rect 1788 8245 1816 8246
rect 1788 8219 1789 8245
rect 1789 8219 1815 8245
rect 1815 8219 1816 8245
rect 1788 8218 1816 8219
rect 854 8078 882 8106
rect 1246 8105 1274 8106
rect 1246 8079 1247 8105
rect 1247 8079 1273 8105
rect 1273 8079 1274 8105
rect 1246 8078 1274 8079
rect 1022 7937 1050 7938
rect 1022 7911 1023 7937
rect 1023 7911 1049 7937
rect 1049 7911 1050 7937
rect 1022 7910 1050 7911
rect 1862 7910 1890 7938
rect 1684 7461 1712 7462
rect 1684 7435 1685 7461
rect 1685 7435 1711 7461
rect 1711 7435 1712 7461
rect 1684 7434 1712 7435
rect 1736 7461 1764 7462
rect 1736 7435 1737 7461
rect 1737 7435 1763 7461
rect 1763 7435 1764 7461
rect 1736 7434 1764 7435
rect 1788 7461 1816 7462
rect 1788 7435 1789 7461
rect 1789 7435 1815 7461
rect 1815 7435 1816 7461
rect 1788 7434 1816 7435
rect 1684 6677 1712 6678
rect 1684 6651 1685 6677
rect 1685 6651 1711 6677
rect 1711 6651 1712 6677
rect 1684 6650 1712 6651
rect 1736 6677 1764 6678
rect 1736 6651 1737 6677
rect 1737 6651 1763 6677
rect 1763 6651 1764 6677
rect 1736 6650 1764 6651
rect 1788 6677 1816 6678
rect 1788 6651 1789 6677
rect 1789 6651 1815 6677
rect 1815 6651 1816 6677
rect 1788 6650 1816 6651
rect 854 6174 882 6202
rect 1246 6174 1274 6202
rect 1684 5893 1712 5894
rect 1684 5867 1685 5893
rect 1685 5867 1711 5893
rect 1711 5867 1712 5893
rect 1684 5866 1712 5867
rect 1736 5893 1764 5894
rect 1736 5867 1737 5893
rect 1737 5867 1763 5893
rect 1763 5867 1764 5893
rect 1736 5866 1764 5867
rect 1788 5893 1816 5894
rect 1788 5867 1789 5893
rect 1789 5867 1815 5893
rect 1815 5867 1816 5893
rect 1788 5866 1816 5867
rect 7406 8358 7434 8386
rect 7910 9198 7938 9226
rect 3840 8245 3868 8246
rect 3840 8219 3841 8245
rect 3841 8219 3867 8245
rect 3867 8219 3868 8245
rect 3840 8218 3868 8219
rect 3892 8245 3920 8246
rect 3892 8219 3893 8245
rect 3893 8219 3919 8245
rect 3919 8219 3920 8245
rect 3892 8218 3920 8219
rect 3944 8245 3972 8246
rect 3944 8219 3945 8245
rect 3945 8219 3971 8245
rect 3971 8219 3972 8245
rect 3944 8218 3972 8219
rect 5996 8245 6024 8246
rect 5996 8219 5997 8245
rect 5997 8219 6023 8245
rect 6023 8219 6024 8245
rect 5996 8218 6024 8219
rect 6048 8245 6076 8246
rect 6048 8219 6049 8245
rect 6049 8219 6075 8245
rect 6075 8219 6076 8245
rect 6048 8218 6076 8219
rect 6100 8245 6128 8246
rect 6100 8219 6101 8245
rect 6101 8219 6127 8245
rect 6127 8219 6128 8245
rect 6100 8218 6128 8219
rect 5446 7966 5474 7994
rect 2762 7853 2790 7854
rect 2762 7827 2763 7853
rect 2763 7827 2789 7853
rect 2789 7827 2790 7853
rect 2762 7826 2790 7827
rect 2814 7853 2842 7854
rect 2814 7827 2815 7853
rect 2815 7827 2841 7853
rect 2841 7827 2842 7853
rect 2814 7826 2842 7827
rect 2866 7853 2894 7854
rect 2866 7827 2867 7853
rect 2867 7827 2893 7853
rect 2893 7827 2894 7853
rect 2866 7826 2894 7827
rect 4918 7853 4946 7854
rect 4918 7827 4919 7853
rect 4919 7827 4945 7853
rect 4945 7827 4946 7853
rect 4918 7826 4946 7827
rect 4970 7853 4998 7854
rect 4970 7827 4971 7853
rect 4971 7827 4997 7853
rect 4997 7827 4998 7853
rect 4970 7826 4998 7827
rect 5022 7853 5050 7854
rect 5022 7827 5023 7853
rect 5023 7827 5049 7853
rect 5049 7827 5050 7853
rect 5022 7826 5050 7827
rect 3430 7657 3458 7658
rect 3430 7631 3431 7657
rect 3431 7631 3457 7657
rect 3457 7631 3458 7657
rect 3430 7630 3458 7631
rect 3840 7461 3868 7462
rect 3840 7435 3841 7461
rect 3841 7435 3867 7461
rect 3867 7435 3868 7461
rect 3840 7434 3868 7435
rect 3892 7461 3920 7462
rect 3892 7435 3893 7461
rect 3893 7435 3919 7461
rect 3919 7435 3920 7461
rect 3892 7434 3920 7435
rect 3944 7461 3972 7462
rect 3944 7435 3945 7461
rect 3945 7435 3971 7461
rect 3971 7435 3972 7461
rect 4494 7462 4522 7490
rect 3944 7434 3972 7435
rect 3094 7350 3122 7378
rect 3598 7350 3626 7378
rect 3374 7126 3402 7154
rect 2762 7069 2790 7070
rect 2762 7043 2763 7069
rect 2763 7043 2789 7069
rect 2789 7043 2790 7069
rect 2762 7042 2790 7043
rect 2814 7069 2842 7070
rect 2814 7043 2815 7069
rect 2815 7043 2841 7069
rect 2841 7043 2842 7069
rect 2814 7042 2842 7043
rect 2866 7069 2894 7070
rect 2866 7043 2867 7069
rect 2867 7043 2893 7069
rect 2893 7043 2894 7069
rect 2866 7042 2894 7043
rect 2478 6174 2506 6202
rect 1974 6089 2002 6090
rect 1974 6063 1975 6089
rect 1975 6063 2001 6089
rect 2001 6063 2002 6089
rect 1974 6062 2002 6063
rect 2982 6817 3010 6818
rect 2982 6791 2983 6817
rect 2983 6791 3009 6817
rect 3009 6791 3010 6817
rect 2982 6790 3010 6791
rect 2762 6285 2790 6286
rect 2762 6259 2763 6285
rect 2763 6259 2789 6285
rect 2789 6259 2790 6285
rect 2762 6258 2790 6259
rect 2814 6285 2842 6286
rect 2814 6259 2815 6285
rect 2815 6259 2841 6285
rect 2841 6259 2842 6285
rect 2814 6258 2842 6259
rect 2866 6285 2894 6286
rect 2866 6259 2867 6285
rect 2867 6259 2893 6285
rect 2893 6259 2894 6285
rect 2866 6258 2894 6259
rect 2702 6062 2730 6090
rect 2310 5950 2338 5978
rect 4942 7574 4970 7602
rect 4326 7350 4354 7378
rect 4774 7462 4802 7490
rect 3934 7153 3962 7154
rect 3934 7127 3935 7153
rect 3935 7127 3961 7153
rect 3961 7127 3962 7153
rect 3934 7126 3962 7127
rect 4046 6734 4074 6762
rect 3840 6677 3868 6678
rect 3840 6651 3841 6677
rect 3841 6651 3867 6677
rect 3867 6651 3868 6677
rect 3840 6650 3868 6651
rect 3892 6677 3920 6678
rect 3892 6651 3893 6677
rect 3893 6651 3919 6677
rect 3919 6651 3920 6677
rect 3892 6650 3920 6651
rect 3944 6677 3972 6678
rect 3944 6651 3945 6677
rect 3945 6651 3971 6677
rect 3971 6651 3972 6677
rect 3944 6650 3972 6651
rect 4214 6481 4242 6482
rect 4214 6455 4215 6481
rect 4215 6455 4241 6481
rect 4241 6455 4242 6481
rect 4214 6454 4242 6455
rect 4046 6398 4074 6426
rect 1022 3793 1050 3794
rect 1022 3767 1023 3793
rect 1023 3767 1049 3793
rect 1049 3767 1050 3793
rect 1022 3766 1050 3767
rect 910 3710 938 3738
rect 1078 3737 1106 3738
rect 1078 3711 1079 3737
rect 1079 3711 1105 3737
rect 1105 3711 1106 3737
rect 1078 3710 1106 3711
rect 1638 5446 1666 5474
rect 2762 5501 2790 5502
rect 2762 5475 2763 5501
rect 2763 5475 2789 5501
rect 2789 5475 2790 5501
rect 2762 5474 2790 5475
rect 2814 5501 2842 5502
rect 2814 5475 2815 5501
rect 2815 5475 2841 5501
rect 2841 5475 2842 5501
rect 2814 5474 2842 5475
rect 2866 5501 2894 5502
rect 2866 5475 2867 5501
rect 2867 5475 2893 5501
rect 2893 5475 2894 5501
rect 2866 5474 2894 5475
rect 2590 5278 2618 5306
rect 1684 5109 1712 5110
rect 1684 5083 1685 5109
rect 1685 5083 1711 5109
rect 1711 5083 1712 5109
rect 1684 5082 1712 5083
rect 1736 5109 1764 5110
rect 1736 5083 1737 5109
rect 1737 5083 1763 5109
rect 1763 5083 1764 5109
rect 1736 5082 1764 5083
rect 1788 5109 1816 5110
rect 1788 5083 1789 5109
rect 1789 5083 1815 5109
rect 1815 5083 1816 5109
rect 1788 5082 1816 5083
rect 1684 4325 1712 4326
rect 1684 4299 1685 4325
rect 1685 4299 1711 4325
rect 1711 4299 1712 4325
rect 1684 4298 1712 4299
rect 1736 4325 1764 4326
rect 1736 4299 1737 4325
rect 1737 4299 1763 4325
rect 1763 4299 1764 4325
rect 1736 4298 1764 4299
rect 1788 4325 1816 4326
rect 1788 4299 1789 4325
rect 1789 4299 1815 4325
rect 1815 4299 1816 4325
rect 1788 4298 1816 4299
rect 1750 4046 1778 4074
rect 1302 3766 1330 3794
rect 1414 3654 1442 3682
rect 2142 4550 2170 4578
rect 1862 4073 1890 4074
rect 1862 4047 1863 4073
rect 1863 4047 1889 4073
rect 1889 4047 1890 4073
rect 1862 4046 1890 4047
rect 2534 4550 2562 4578
rect 2702 4998 2730 5026
rect 2870 5249 2898 5250
rect 2870 5223 2871 5249
rect 2871 5223 2897 5249
rect 2897 5223 2898 5249
rect 2870 5222 2898 5223
rect 2982 4998 3010 5026
rect 3094 5054 3122 5082
rect 3038 4942 3066 4970
rect 2762 4717 2790 4718
rect 2762 4691 2763 4717
rect 2763 4691 2789 4717
rect 2789 4691 2790 4717
rect 2762 4690 2790 4691
rect 2814 4717 2842 4718
rect 2814 4691 2815 4717
rect 2815 4691 2841 4717
rect 2841 4691 2842 4717
rect 2814 4690 2842 4691
rect 2866 4717 2894 4718
rect 2866 4691 2867 4717
rect 2867 4691 2893 4717
rect 2893 4691 2894 4717
rect 2866 4690 2894 4691
rect 2758 4577 2786 4578
rect 2758 4551 2759 4577
rect 2759 4551 2785 4577
rect 2785 4551 2786 4577
rect 2758 4550 2786 4551
rect 1862 3766 1890 3794
rect 2478 3793 2506 3794
rect 2478 3767 2479 3793
rect 2479 3767 2505 3793
rect 2505 3767 2506 3793
rect 2478 3766 2506 3767
rect 1750 3654 1778 3682
rect 1684 3541 1712 3542
rect 1684 3515 1685 3541
rect 1685 3515 1711 3541
rect 1711 3515 1712 3541
rect 1684 3514 1712 3515
rect 1736 3541 1764 3542
rect 1736 3515 1737 3541
rect 1737 3515 1763 3541
rect 1763 3515 1764 3541
rect 1736 3514 1764 3515
rect 1788 3541 1816 3542
rect 1788 3515 1789 3541
rect 1789 3515 1815 3541
rect 1815 3515 1816 3541
rect 1788 3514 1816 3515
rect 2030 3486 2058 3514
rect 2310 3737 2338 3738
rect 2310 3711 2311 3737
rect 2311 3711 2337 3737
rect 2337 3711 2338 3737
rect 2310 3710 2338 3711
rect 2198 3654 2226 3682
rect 2198 3430 2226 3458
rect 1526 3374 1554 3402
rect 1302 3262 1330 3290
rect 2534 3486 2562 3514
rect 2870 4494 2898 4522
rect 2254 3374 2282 3402
rect 1918 3262 1946 3290
rect 1134 2953 1162 2954
rect 1134 2927 1135 2953
rect 1135 2927 1161 2953
rect 1161 2927 1162 2953
rect 1134 2926 1162 2927
rect 1684 2757 1712 2758
rect 1684 2731 1685 2757
rect 1685 2731 1711 2757
rect 1711 2731 1712 2757
rect 1684 2730 1712 2731
rect 1736 2757 1764 2758
rect 1736 2731 1737 2757
rect 1737 2731 1763 2757
rect 1763 2731 1764 2757
rect 1736 2730 1764 2731
rect 1788 2757 1816 2758
rect 1788 2731 1789 2757
rect 1789 2731 1815 2757
rect 1815 2731 1816 2757
rect 1788 2730 1816 2731
rect 1684 1973 1712 1974
rect 1684 1947 1685 1973
rect 1685 1947 1711 1973
rect 1711 1947 1712 1973
rect 1684 1946 1712 1947
rect 1736 1973 1764 1974
rect 1736 1947 1737 1973
rect 1737 1947 1763 1973
rect 1763 1947 1764 1973
rect 1736 1946 1764 1947
rect 1788 1973 1816 1974
rect 1788 1947 1789 1973
rect 1789 1947 1815 1973
rect 1815 1947 1816 1973
rect 1788 1946 1816 1947
rect 2762 3933 2790 3934
rect 2762 3907 2763 3933
rect 2763 3907 2789 3933
rect 2789 3907 2790 3933
rect 2762 3906 2790 3907
rect 2814 3933 2842 3934
rect 2814 3907 2815 3933
rect 2815 3907 2841 3933
rect 2841 3907 2842 3933
rect 2814 3906 2842 3907
rect 2866 3933 2894 3934
rect 2866 3907 2867 3933
rect 2867 3907 2893 3933
rect 2893 3907 2894 3933
rect 2866 3906 2894 3907
rect 2762 3149 2790 3150
rect 2762 3123 2763 3149
rect 2763 3123 2789 3149
rect 2789 3123 2790 3149
rect 2762 3122 2790 3123
rect 2814 3149 2842 3150
rect 2814 3123 2815 3149
rect 2815 3123 2841 3149
rect 2841 3123 2842 3149
rect 2814 3122 2842 3123
rect 2866 3149 2894 3150
rect 2866 3123 2867 3149
rect 2867 3123 2893 3149
rect 2893 3123 2894 3149
rect 2866 3122 2894 3123
rect 2702 3038 2730 3066
rect 3038 4521 3066 4522
rect 3038 4495 3039 4521
rect 3039 4495 3065 4521
rect 3065 4495 3066 4521
rect 3038 4494 3066 4495
rect 2982 3822 3010 3850
rect 3206 4606 3234 4634
rect 3318 5390 3346 5418
rect 3486 5305 3514 5306
rect 3486 5279 3487 5305
rect 3487 5279 3513 5305
rect 3513 5279 3514 5305
rect 3486 5278 3514 5279
rect 3598 5305 3626 5306
rect 3598 5279 3599 5305
rect 3599 5279 3625 5305
rect 3625 5279 3626 5305
rect 3598 5278 3626 5279
rect 3318 5054 3346 5082
rect 4270 6398 4298 6426
rect 4662 7182 4690 7210
rect 4494 6929 4522 6930
rect 4494 6903 4495 6929
rect 4495 6903 4521 6929
rect 4521 6903 4522 6929
rect 4494 6902 4522 6903
rect 6118 7993 6146 7994
rect 6118 7967 6119 7993
rect 6119 7967 6145 7993
rect 6145 7967 6146 7993
rect 6118 7966 6146 7967
rect 7406 7993 7434 7994
rect 7406 7967 7407 7993
rect 7407 7967 7433 7993
rect 7433 7967 7434 7993
rect 7406 7966 7434 7967
rect 5446 7601 5474 7602
rect 5446 7575 5447 7601
rect 5447 7575 5473 7601
rect 5473 7575 5474 7601
rect 5446 7574 5474 7575
rect 5782 7630 5810 7658
rect 4998 7462 5026 7490
rect 4774 7126 4802 7154
rect 4918 7069 4946 7070
rect 4918 7043 4919 7069
rect 4919 7043 4945 7069
rect 4945 7043 4946 7069
rect 4918 7042 4946 7043
rect 4970 7069 4998 7070
rect 4970 7043 4971 7069
rect 4971 7043 4997 7069
rect 4997 7043 4998 7069
rect 4970 7042 4998 7043
rect 5022 7069 5050 7070
rect 5022 7043 5023 7069
rect 5023 7043 5049 7069
rect 5049 7043 5050 7069
rect 5022 7042 5050 7043
rect 5278 7238 5306 7266
rect 5166 7153 5194 7154
rect 5166 7127 5167 7153
rect 5167 7127 5193 7153
rect 5193 7127 5194 7153
rect 5166 7126 5194 7127
rect 4998 6958 5026 6986
rect 4438 6734 4466 6762
rect 4718 6734 4746 6762
rect 4662 6566 4690 6594
rect 4382 6510 4410 6538
rect 4606 6510 4634 6538
rect 3990 6089 4018 6090
rect 3990 6063 3991 6089
rect 3991 6063 4017 6089
rect 4017 6063 4018 6089
rect 3990 6062 4018 6063
rect 3840 5893 3868 5894
rect 3840 5867 3841 5893
rect 3841 5867 3867 5893
rect 3867 5867 3868 5893
rect 3840 5866 3868 5867
rect 3892 5893 3920 5894
rect 3892 5867 3893 5893
rect 3893 5867 3919 5893
rect 3919 5867 3920 5893
rect 3892 5866 3920 5867
rect 3944 5893 3972 5894
rect 3944 5867 3945 5893
rect 3945 5867 3971 5893
rect 3971 5867 3972 5893
rect 3944 5866 3972 5867
rect 3710 5249 3738 5250
rect 3710 5223 3711 5249
rect 3711 5223 3737 5249
rect 3737 5223 3738 5249
rect 3710 5222 3738 5223
rect 3654 4969 3682 4970
rect 3654 4943 3655 4969
rect 3655 4943 3681 4969
rect 3681 4943 3682 4969
rect 3654 4942 3682 4943
rect 3710 4606 3738 4634
rect 3934 5222 3962 5250
rect 4046 5166 4074 5194
rect 4606 6425 4634 6426
rect 4606 6399 4607 6425
rect 4607 6399 4633 6425
rect 4633 6399 4634 6425
rect 4606 6398 4634 6399
rect 4326 6118 4354 6146
rect 4382 6089 4410 6090
rect 4382 6063 4383 6089
rect 4383 6063 4409 6089
rect 4409 6063 4410 6089
rect 4382 6062 4410 6063
rect 4102 5222 4130 5250
rect 5166 6902 5194 6930
rect 5110 6761 5138 6762
rect 5110 6735 5111 6761
rect 5111 6735 5137 6761
rect 5137 6735 5138 6761
rect 5110 6734 5138 6735
rect 5558 7209 5586 7210
rect 5558 7183 5559 7209
rect 5559 7183 5585 7209
rect 5585 7183 5586 7209
rect 5558 7182 5586 7183
rect 5670 7153 5698 7154
rect 5670 7127 5671 7153
rect 5671 7127 5697 7153
rect 5697 7127 5698 7153
rect 5670 7126 5698 7127
rect 5222 6790 5250 6818
rect 4918 6285 4946 6286
rect 4918 6259 4919 6285
rect 4919 6259 4945 6285
rect 4945 6259 4946 6285
rect 4918 6258 4946 6259
rect 4970 6285 4998 6286
rect 4970 6259 4971 6285
rect 4971 6259 4997 6285
rect 4997 6259 4998 6285
rect 4970 6258 4998 6259
rect 5022 6285 5050 6286
rect 5022 6259 5023 6285
rect 5023 6259 5049 6285
rect 5049 6259 5050 6285
rect 5022 6258 5050 6259
rect 5166 6230 5194 6258
rect 4830 6201 4858 6202
rect 4830 6175 4831 6201
rect 4831 6175 4857 6201
rect 4857 6175 4858 6201
rect 4830 6174 4858 6175
rect 5054 6174 5082 6202
rect 4662 6118 4690 6146
rect 4550 5670 4578 5698
rect 4438 5334 4466 5362
rect 4270 5222 4298 5250
rect 3840 5109 3868 5110
rect 3840 5083 3841 5109
rect 3841 5083 3867 5109
rect 3867 5083 3868 5109
rect 3840 5082 3868 5083
rect 3892 5109 3920 5110
rect 3892 5083 3893 5109
rect 3893 5083 3919 5109
rect 3919 5083 3920 5109
rect 3892 5082 3920 5083
rect 3944 5109 3972 5110
rect 3944 5083 3945 5109
rect 3945 5083 3971 5109
rect 3971 5083 3972 5109
rect 3944 5082 3972 5083
rect 4102 5054 4130 5082
rect 3840 4325 3868 4326
rect 3840 4299 3841 4325
rect 3841 4299 3867 4325
rect 3867 4299 3868 4325
rect 3840 4298 3868 4299
rect 3892 4325 3920 4326
rect 3892 4299 3893 4325
rect 3893 4299 3919 4325
rect 3919 4299 3920 4325
rect 3892 4298 3920 4299
rect 3944 4325 3972 4326
rect 3944 4299 3945 4325
rect 3945 4299 3971 4325
rect 3971 4299 3972 4325
rect 3944 4298 3972 4299
rect 3094 3766 3122 3794
rect 3150 3737 3178 3738
rect 3150 3711 3151 3737
rect 3151 3711 3177 3737
rect 3177 3711 3178 3737
rect 3150 3710 3178 3711
rect 2142 2926 2170 2954
rect 2814 2926 2842 2954
rect 3038 3486 3066 3514
rect 3094 3457 3122 3458
rect 3094 3431 3095 3457
rect 3095 3431 3121 3457
rect 3121 3431 3122 3457
rect 3094 3430 3122 3431
rect 3094 3065 3122 3066
rect 3094 3039 3095 3065
rect 3095 3039 3121 3065
rect 3121 3039 3122 3065
rect 3094 3038 3122 3039
rect 2478 2590 2506 2618
rect 2926 2617 2954 2618
rect 2926 2591 2927 2617
rect 2927 2591 2953 2617
rect 2953 2591 2954 2617
rect 2926 2590 2954 2591
rect 2590 2561 2618 2562
rect 2590 2535 2591 2561
rect 2591 2535 2617 2561
rect 2617 2535 2618 2561
rect 2590 2534 2618 2535
rect 2982 2534 3010 2562
rect 2762 2365 2790 2366
rect 2762 2339 2763 2365
rect 2763 2339 2789 2365
rect 2789 2339 2790 2365
rect 2762 2338 2790 2339
rect 2814 2365 2842 2366
rect 2814 2339 2815 2365
rect 2815 2339 2841 2365
rect 2841 2339 2842 2365
rect 2814 2338 2842 2339
rect 2866 2365 2894 2366
rect 2866 2339 2867 2365
rect 2867 2339 2893 2365
rect 2893 2339 2894 2365
rect 2866 2338 2894 2339
rect 3206 2870 3234 2898
rect 3654 3710 3682 3738
rect 3878 4017 3906 4018
rect 3878 3991 3879 4017
rect 3879 3991 3905 4017
rect 3905 3991 3906 4017
rect 3878 3990 3906 3991
rect 4550 5278 4578 5306
rect 4494 4046 4522 4074
rect 4550 4942 4578 4970
rect 4942 5950 4970 5978
rect 4886 5697 4914 5698
rect 4886 5671 4887 5697
rect 4887 5671 4913 5697
rect 4913 5671 4914 5697
rect 4886 5670 4914 5671
rect 4998 5697 5026 5698
rect 4998 5671 4999 5697
rect 4999 5671 5025 5697
rect 5025 5671 5026 5697
rect 4998 5670 5026 5671
rect 5334 6622 5362 6650
rect 5278 6566 5306 6594
rect 5334 6537 5362 6538
rect 5334 6511 5335 6537
rect 5335 6511 5361 6537
rect 5361 6511 5362 6537
rect 5334 6510 5362 6511
rect 5278 6398 5306 6426
rect 5502 6510 5530 6538
rect 5278 6286 5306 6314
rect 5390 6174 5418 6202
rect 5166 5809 5194 5810
rect 5166 5783 5167 5809
rect 5167 5783 5193 5809
rect 5193 5783 5194 5809
rect 5166 5782 5194 5783
rect 5110 5670 5138 5698
rect 4918 5501 4946 5502
rect 4918 5475 4919 5501
rect 4919 5475 4945 5501
rect 4945 5475 4946 5501
rect 4918 5474 4946 5475
rect 4970 5501 4998 5502
rect 4970 5475 4971 5501
rect 4971 5475 4997 5501
rect 4997 5475 4998 5501
rect 4970 5474 4998 5475
rect 5022 5501 5050 5502
rect 5022 5475 5023 5501
rect 5023 5475 5049 5501
rect 5049 5475 5050 5501
rect 5022 5474 5050 5475
rect 4774 5361 4802 5362
rect 4774 5335 4775 5361
rect 4775 5335 4801 5361
rect 4801 5335 4802 5361
rect 4774 5334 4802 5335
rect 4830 5278 4858 5306
rect 4774 5166 4802 5194
rect 4942 5305 4970 5306
rect 4942 5279 4943 5305
rect 4943 5279 4969 5305
rect 4969 5279 4970 5305
rect 4942 5278 4970 5279
rect 5166 5558 5194 5586
rect 5278 5977 5306 5978
rect 5278 5951 5279 5977
rect 5279 5951 5305 5977
rect 5305 5951 5306 5977
rect 5278 5950 5306 5951
rect 5334 5446 5362 5474
rect 5222 5278 5250 5306
rect 5334 5334 5362 5362
rect 4918 4717 4946 4718
rect 4918 4691 4919 4717
rect 4919 4691 4945 4717
rect 4945 4691 4946 4717
rect 4918 4690 4946 4691
rect 4970 4717 4998 4718
rect 4970 4691 4971 4717
rect 4971 4691 4997 4717
rect 4997 4691 4998 4717
rect 4970 4690 4998 4691
rect 5022 4717 5050 4718
rect 5022 4691 5023 4717
rect 5023 4691 5049 4717
rect 5049 4691 5050 4717
rect 5022 4690 5050 4691
rect 5558 6286 5586 6314
rect 6230 7574 6258 7602
rect 5996 7461 6024 7462
rect 5996 7435 5997 7461
rect 5997 7435 6023 7461
rect 6023 7435 6024 7461
rect 5996 7434 6024 7435
rect 6048 7461 6076 7462
rect 6048 7435 6049 7461
rect 6049 7435 6075 7461
rect 6075 7435 6076 7461
rect 6048 7434 6076 7435
rect 6100 7461 6128 7462
rect 6100 7435 6101 7461
rect 6101 7435 6127 7461
rect 6127 7435 6128 7461
rect 6100 7434 6128 7435
rect 5894 7265 5922 7266
rect 5894 7239 5895 7265
rect 5895 7239 5921 7265
rect 5921 7239 5922 7265
rect 5894 7238 5922 7239
rect 5838 7126 5866 7154
rect 7074 7853 7102 7854
rect 7074 7827 7075 7853
rect 7075 7827 7101 7853
rect 7101 7827 7102 7853
rect 7074 7826 7102 7827
rect 7126 7853 7154 7854
rect 7126 7827 7127 7853
rect 7127 7827 7153 7853
rect 7153 7827 7154 7853
rect 7126 7826 7154 7827
rect 7178 7853 7206 7854
rect 7178 7827 7179 7853
rect 7179 7827 7205 7853
rect 7205 7827 7206 7853
rect 7178 7826 7206 7827
rect 8582 8358 8610 8386
rect 8152 8245 8180 8246
rect 8152 8219 8153 8245
rect 8153 8219 8179 8245
rect 8179 8219 8180 8245
rect 8152 8218 8180 8219
rect 8204 8245 8232 8246
rect 8204 8219 8205 8245
rect 8205 8219 8231 8245
rect 8231 8219 8232 8245
rect 8204 8218 8232 8219
rect 8256 8245 8284 8246
rect 8256 8219 8257 8245
rect 8257 8219 8283 8245
rect 8283 8219 8284 8245
rect 8256 8218 8284 8219
rect 8582 8078 8610 8106
rect 8190 8049 8218 8050
rect 8190 8023 8191 8049
rect 8191 8023 8217 8049
rect 8217 8023 8218 8049
rect 8190 8022 8218 8023
rect 8862 8105 8890 8106
rect 8862 8079 8863 8105
rect 8863 8079 8889 8105
rect 8889 8079 8890 8105
rect 8862 8078 8890 8079
rect 8806 8022 8834 8050
rect 6902 7657 6930 7658
rect 6902 7631 6903 7657
rect 6903 7631 6929 7657
rect 6929 7631 6930 7657
rect 6902 7630 6930 7631
rect 7574 7630 7602 7658
rect 6510 7601 6538 7602
rect 6510 7575 6511 7601
rect 6511 7575 6537 7601
rect 6537 7575 6538 7601
rect 6510 7574 6538 7575
rect 6398 7238 6426 7266
rect 6006 7153 6034 7154
rect 6006 7127 6007 7153
rect 6007 7127 6033 7153
rect 6033 7127 6034 7153
rect 6006 7126 6034 7127
rect 5838 6958 5866 6986
rect 5670 6342 5698 6370
rect 7238 7265 7266 7266
rect 7238 7239 7239 7265
rect 7239 7239 7265 7265
rect 7265 7239 7266 7265
rect 7238 7238 7266 7239
rect 5782 6678 5810 6706
rect 5950 6873 5978 6874
rect 5950 6847 5951 6873
rect 5951 6847 5977 6873
rect 5977 6847 5978 6873
rect 5950 6846 5978 6847
rect 6062 6761 6090 6762
rect 6062 6735 6063 6761
rect 6063 6735 6089 6761
rect 6089 6735 6090 6761
rect 6062 6734 6090 6735
rect 6174 6873 6202 6874
rect 6174 6847 6175 6873
rect 6175 6847 6201 6873
rect 6201 6847 6202 6873
rect 6174 6846 6202 6847
rect 5996 6677 6024 6678
rect 5996 6651 5997 6677
rect 5997 6651 6023 6677
rect 6023 6651 6024 6677
rect 5996 6650 6024 6651
rect 6048 6677 6076 6678
rect 6048 6651 6049 6677
rect 6049 6651 6075 6677
rect 6075 6651 6076 6677
rect 6048 6650 6076 6651
rect 6100 6677 6128 6678
rect 6100 6651 6101 6677
rect 6101 6651 6127 6677
rect 6127 6651 6128 6677
rect 6100 6650 6128 6651
rect 6174 6566 6202 6594
rect 6454 7209 6482 7210
rect 6454 7183 6455 7209
rect 6455 7183 6481 7209
rect 6481 7183 6482 7209
rect 6454 7182 6482 7183
rect 6678 7126 6706 7154
rect 6006 6481 6034 6482
rect 6006 6455 6007 6481
rect 6007 6455 6033 6481
rect 6033 6455 6034 6481
rect 6006 6454 6034 6455
rect 5838 6230 5866 6258
rect 5950 6062 5978 6090
rect 5726 6006 5754 6034
rect 5894 5977 5922 5978
rect 5894 5951 5895 5977
rect 5895 5951 5921 5977
rect 5921 5951 5922 5977
rect 5894 5950 5922 5951
rect 6174 6425 6202 6426
rect 6174 6399 6175 6425
rect 6175 6399 6201 6425
rect 6201 6399 6202 6425
rect 6174 6398 6202 6399
rect 6006 5950 6034 5978
rect 6062 6286 6090 6314
rect 6510 6846 6538 6874
rect 7126 7209 7154 7210
rect 7126 7183 7127 7209
rect 7127 7183 7153 7209
rect 7153 7183 7154 7209
rect 7126 7182 7154 7183
rect 7074 7069 7102 7070
rect 7074 7043 7075 7069
rect 7075 7043 7101 7069
rect 7101 7043 7102 7069
rect 7074 7042 7102 7043
rect 7126 7069 7154 7070
rect 7126 7043 7127 7069
rect 7127 7043 7153 7069
rect 7153 7043 7154 7069
rect 7126 7042 7154 7043
rect 7178 7069 7206 7070
rect 7178 7043 7179 7069
rect 7179 7043 7205 7069
rect 7205 7043 7206 7069
rect 7178 7042 7206 7043
rect 6566 6566 6594 6594
rect 6062 6006 6090 6034
rect 5996 5893 6024 5894
rect 5996 5867 5997 5893
rect 5997 5867 6023 5893
rect 6023 5867 6024 5893
rect 5996 5866 6024 5867
rect 6048 5893 6076 5894
rect 6048 5867 6049 5893
rect 6049 5867 6075 5893
rect 6075 5867 6076 5893
rect 6048 5866 6076 5867
rect 6100 5893 6128 5894
rect 6100 5867 6101 5893
rect 6101 5867 6127 5893
rect 6127 5867 6128 5893
rect 6100 5866 6128 5867
rect 5446 5222 5474 5250
rect 4438 3990 4466 4018
rect 3822 3710 3850 3738
rect 3318 2646 3346 2674
rect 3840 3541 3868 3542
rect 3840 3515 3841 3541
rect 3841 3515 3867 3541
rect 3867 3515 3868 3541
rect 3840 3514 3868 3515
rect 3892 3541 3920 3542
rect 3892 3515 3893 3541
rect 3893 3515 3919 3541
rect 3919 3515 3920 3541
rect 3892 3514 3920 3515
rect 3944 3541 3972 3542
rect 3944 3515 3945 3541
rect 3945 3515 3971 3541
rect 3971 3515 3972 3541
rect 3944 3514 3972 3515
rect 3654 3345 3682 3346
rect 3654 3319 3655 3345
rect 3655 3319 3681 3345
rect 3681 3319 3682 3345
rect 3654 3318 3682 3319
rect 3486 3065 3514 3066
rect 3486 3039 3487 3065
rect 3487 3039 3513 3065
rect 3513 3039 3514 3065
rect 3486 3038 3514 3039
rect 3710 2926 3738 2954
rect 3094 2142 3122 2170
rect 3766 2870 3794 2898
rect 3934 3318 3962 3346
rect 4214 3262 4242 3290
rect 4270 3094 4298 3122
rect 4942 4073 4970 4074
rect 4942 4047 4943 4073
rect 4943 4047 4969 4073
rect 4969 4047 4970 4073
rect 4942 4046 4970 4047
rect 5390 4465 5418 4466
rect 5390 4439 5391 4465
rect 5391 4439 5417 4465
rect 5417 4439 5418 4465
rect 5390 4438 5418 4439
rect 5222 3990 5250 4018
rect 4918 3933 4946 3934
rect 4918 3907 4919 3933
rect 4919 3907 4945 3933
rect 4945 3907 4946 3933
rect 4918 3906 4946 3907
rect 4970 3933 4998 3934
rect 4970 3907 4971 3933
rect 4971 3907 4997 3933
rect 4997 3907 4998 3933
rect 4970 3906 4998 3907
rect 5022 3933 5050 3934
rect 5022 3907 5023 3933
rect 5023 3907 5049 3933
rect 5049 3907 5050 3933
rect 5022 3906 5050 3907
rect 6286 5782 6314 5810
rect 5950 5670 5978 5698
rect 5670 5585 5698 5586
rect 5670 5559 5671 5585
rect 5671 5559 5697 5585
rect 5697 5559 5698 5585
rect 5670 5558 5698 5559
rect 6958 6622 6986 6650
rect 8414 7657 8442 7658
rect 8414 7631 8415 7657
rect 8415 7631 8441 7657
rect 8441 7631 8442 7657
rect 8414 7630 8442 7631
rect 8152 7461 8180 7462
rect 8152 7435 8153 7461
rect 8153 7435 8179 7461
rect 8179 7435 8180 7461
rect 8152 7434 8180 7435
rect 8204 7461 8232 7462
rect 8204 7435 8205 7461
rect 8205 7435 8231 7461
rect 8231 7435 8232 7461
rect 8204 7434 8232 7435
rect 8256 7461 8284 7462
rect 8256 7435 8257 7461
rect 8257 7435 8283 7461
rect 8283 7435 8284 7461
rect 8256 7434 8284 7435
rect 7518 7182 7546 7210
rect 7294 6622 7322 6650
rect 6958 6342 6986 6370
rect 7014 6481 7042 6482
rect 7014 6455 7015 6481
rect 7015 6455 7041 6481
rect 7041 6455 7042 6481
rect 7014 6454 7042 6455
rect 6566 6062 6594 6090
rect 5614 5334 5642 5362
rect 5950 5502 5978 5530
rect 5726 4998 5754 5026
rect 6174 5558 6202 5586
rect 6230 5502 6258 5530
rect 5996 5109 6024 5110
rect 5996 5083 5997 5109
rect 5997 5083 6023 5109
rect 6023 5083 6024 5109
rect 5996 5082 6024 5083
rect 6048 5109 6076 5110
rect 6048 5083 6049 5109
rect 6049 5083 6075 5109
rect 6075 5083 6076 5109
rect 6048 5082 6076 5083
rect 6100 5109 6128 5110
rect 6100 5083 6101 5109
rect 6101 5083 6127 5109
rect 6127 5083 6128 5109
rect 6100 5082 6128 5083
rect 6174 4998 6202 5026
rect 6118 4942 6146 4970
rect 5894 4438 5922 4466
rect 5996 4325 6024 4326
rect 5996 4299 5997 4325
rect 5997 4299 6023 4325
rect 6023 4299 6024 4325
rect 5996 4298 6024 4299
rect 6048 4325 6076 4326
rect 6048 4299 6049 4325
rect 6049 4299 6075 4325
rect 6075 4299 6076 4325
rect 6048 4298 6076 4299
rect 6100 4325 6128 4326
rect 6100 4299 6101 4325
rect 6101 4299 6127 4325
rect 6127 4299 6128 4325
rect 6100 4298 6128 4299
rect 6006 4102 6034 4130
rect 5502 4046 5530 4074
rect 5894 3990 5922 4018
rect 6902 6118 6930 6146
rect 7294 6425 7322 6426
rect 7294 6399 7295 6425
rect 7295 6399 7321 6425
rect 7321 6399 7322 6425
rect 7294 6398 7322 6399
rect 7126 6369 7154 6370
rect 7126 6343 7127 6369
rect 7127 6343 7153 6369
rect 7153 6343 7154 6369
rect 7126 6342 7154 6343
rect 7074 6285 7102 6286
rect 7074 6259 7075 6285
rect 7075 6259 7101 6285
rect 7101 6259 7102 6285
rect 7074 6258 7102 6259
rect 7126 6285 7154 6286
rect 7126 6259 7127 6285
rect 7127 6259 7153 6285
rect 7153 6259 7154 6285
rect 7126 6258 7154 6259
rect 7178 6285 7206 6286
rect 7178 6259 7179 6285
rect 7179 6259 7205 6285
rect 7205 6259 7206 6285
rect 7178 6258 7206 6259
rect 6734 5641 6762 5642
rect 6734 5615 6735 5641
rect 6735 5615 6761 5641
rect 6761 5615 6762 5641
rect 6734 5614 6762 5615
rect 6342 5558 6370 5586
rect 6734 5390 6762 5418
rect 7182 5838 7210 5866
rect 7070 5641 7098 5642
rect 7070 5615 7071 5641
rect 7071 5615 7097 5641
rect 7097 5615 7098 5641
rect 7070 5614 7098 5615
rect 7074 5501 7102 5502
rect 7074 5475 7075 5501
rect 7075 5475 7101 5501
rect 7101 5475 7102 5501
rect 7074 5474 7102 5475
rect 7126 5501 7154 5502
rect 7126 5475 7127 5501
rect 7127 5475 7153 5501
rect 7153 5475 7154 5501
rect 7126 5474 7154 5475
rect 7178 5501 7206 5502
rect 7178 5475 7179 5501
rect 7179 5475 7205 5501
rect 7205 5475 7206 5501
rect 7178 5474 7206 5475
rect 7182 5390 7210 5418
rect 7406 6510 7434 6538
rect 7350 6230 7378 6258
rect 7294 5753 7322 5754
rect 7294 5727 7295 5753
rect 7295 5727 7321 5753
rect 7321 5727 7322 5753
rect 7294 5726 7322 5727
rect 7406 5614 7434 5642
rect 7966 7209 7994 7210
rect 7966 7183 7967 7209
rect 7967 7183 7993 7209
rect 7993 7183 7994 7209
rect 7966 7182 7994 7183
rect 8414 6873 8442 6874
rect 8414 6847 8415 6873
rect 8415 6847 8441 6873
rect 8441 6847 8442 6873
rect 8414 6846 8442 6847
rect 7910 6761 7938 6762
rect 7910 6735 7911 6761
rect 7911 6735 7937 6761
rect 7937 6735 7938 6761
rect 7910 6734 7938 6735
rect 8152 6677 8180 6678
rect 8152 6651 8153 6677
rect 8153 6651 8179 6677
rect 8179 6651 8180 6677
rect 8152 6650 8180 6651
rect 8204 6677 8232 6678
rect 8204 6651 8205 6677
rect 8205 6651 8231 6677
rect 8231 6651 8232 6677
rect 8204 6650 8232 6651
rect 8256 6677 8284 6678
rect 8256 6651 8257 6677
rect 8257 6651 8283 6677
rect 8283 6651 8284 6677
rect 8256 6650 8284 6651
rect 8022 6537 8050 6538
rect 8022 6511 8023 6537
rect 8023 6511 8049 6537
rect 8049 6511 8050 6537
rect 8022 6510 8050 6511
rect 9230 7853 9258 7854
rect 9230 7827 9231 7853
rect 9231 7827 9257 7853
rect 9257 7827 9258 7853
rect 9230 7826 9258 7827
rect 9282 7853 9310 7854
rect 9282 7827 9283 7853
rect 9283 7827 9309 7853
rect 9309 7827 9310 7853
rect 9282 7826 9310 7827
rect 9334 7853 9362 7854
rect 9334 7827 9335 7853
rect 9335 7827 9361 7853
rect 9361 7827 9362 7853
rect 9334 7826 9362 7827
rect 8470 6454 8498 6482
rect 8750 7238 8778 7266
rect 8694 6398 8722 6426
rect 8638 6118 8666 6146
rect 7966 6062 7994 6090
rect 7462 5278 7490 5306
rect 6286 4102 6314 4130
rect 5278 3374 5306 3402
rect 4158 3038 4186 3066
rect 4998 3289 5026 3290
rect 4998 3263 4999 3289
rect 4999 3263 5025 3289
rect 5025 3263 5026 3289
rect 4998 3262 5026 3263
rect 4918 3149 4946 3150
rect 4918 3123 4919 3149
rect 4919 3123 4945 3149
rect 4945 3123 4946 3149
rect 4918 3122 4946 3123
rect 4970 3149 4998 3150
rect 4970 3123 4971 3149
rect 4971 3123 4997 3149
rect 4997 3123 4998 3149
rect 4970 3122 4998 3123
rect 5022 3149 5050 3150
rect 5022 3123 5023 3149
rect 5023 3123 5049 3149
rect 5049 3123 5050 3149
rect 5022 3122 5050 3123
rect 5222 3065 5250 3066
rect 5222 3039 5223 3065
rect 5223 3039 5249 3065
rect 5249 3039 5250 3065
rect 5222 3038 5250 3039
rect 4382 2982 4410 3010
rect 4998 3009 5026 3010
rect 4998 2983 4999 3009
rect 4999 2983 5025 3009
rect 5025 2983 5026 3009
rect 4998 2982 5026 2983
rect 3990 2870 4018 2898
rect 4046 2814 4074 2842
rect 3840 2757 3868 2758
rect 3840 2731 3841 2757
rect 3841 2731 3867 2757
rect 3867 2731 3868 2757
rect 3840 2730 3868 2731
rect 3892 2757 3920 2758
rect 3892 2731 3893 2757
rect 3893 2731 3919 2757
rect 3919 2731 3920 2757
rect 3892 2730 3920 2731
rect 3944 2757 3972 2758
rect 3944 2731 3945 2757
rect 3945 2731 3971 2757
rect 3971 2731 3972 2757
rect 3944 2730 3972 2731
rect 3878 2646 3906 2674
rect 4886 2841 4914 2842
rect 4886 2815 4887 2841
rect 4887 2815 4913 2841
rect 4913 2815 4914 2841
rect 4886 2814 4914 2815
rect 3934 2169 3962 2170
rect 3934 2143 3935 2169
rect 3935 2143 3961 2169
rect 3961 2143 3962 2169
rect 3934 2142 3962 2143
rect 3840 1973 3868 1974
rect 3840 1947 3841 1973
rect 3841 1947 3867 1973
rect 3867 1947 3868 1973
rect 3840 1946 3868 1947
rect 3892 1973 3920 1974
rect 3892 1947 3893 1973
rect 3893 1947 3919 1973
rect 3919 1947 3920 1973
rect 3892 1946 3920 1947
rect 3944 1973 3972 1974
rect 3944 1947 3945 1973
rect 3945 1947 3971 1973
rect 3971 1947 3972 1973
rect 3944 1946 3972 1947
rect 4326 2561 4354 2562
rect 4326 2535 4327 2561
rect 4327 2535 4353 2561
rect 4353 2535 4354 2561
rect 4326 2534 4354 2535
rect 4718 2449 4746 2450
rect 4718 2423 4719 2449
rect 4719 2423 4745 2449
rect 4745 2423 4746 2449
rect 4718 2422 4746 2423
rect 5996 3541 6024 3542
rect 5996 3515 5997 3541
rect 5997 3515 6023 3541
rect 6023 3515 6024 3541
rect 5996 3514 6024 3515
rect 6048 3541 6076 3542
rect 6048 3515 6049 3541
rect 6049 3515 6075 3541
rect 6075 3515 6076 3541
rect 6048 3514 6076 3515
rect 6100 3541 6128 3542
rect 6100 3515 6101 3541
rect 6101 3515 6127 3541
rect 6127 3515 6128 3541
rect 6100 3514 6128 3515
rect 6062 3401 6090 3402
rect 6062 3375 6063 3401
rect 6063 3375 6089 3401
rect 6089 3375 6090 3401
rect 6062 3374 6090 3375
rect 6230 2870 6258 2898
rect 5996 2757 6024 2758
rect 5996 2731 5997 2757
rect 5997 2731 6023 2757
rect 6023 2731 6024 2757
rect 5996 2730 6024 2731
rect 6048 2757 6076 2758
rect 6048 2731 6049 2757
rect 6049 2731 6075 2757
rect 6075 2731 6076 2757
rect 6048 2730 6076 2731
rect 6100 2757 6128 2758
rect 6100 2731 6101 2757
rect 6101 2731 6127 2757
rect 6127 2731 6128 2757
rect 6100 2730 6128 2731
rect 4998 2590 5026 2618
rect 6006 2617 6034 2618
rect 6006 2591 6007 2617
rect 6007 2591 6033 2617
rect 6033 2591 6034 2617
rect 6006 2590 6034 2591
rect 4918 2365 4946 2366
rect 4918 2339 4919 2365
rect 4919 2339 4945 2365
rect 4945 2339 4946 2365
rect 4918 2338 4946 2339
rect 4970 2365 4998 2366
rect 4970 2339 4971 2365
rect 4971 2339 4997 2365
rect 4997 2339 4998 2365
rect 4970 2338 4998 2339
rect 5022 2365 5050 2366
rect 5022 2339 5023 2365
rect 5023 2339 5049 2365
rect 5049 2339 5050 2365
rect 5022 2338 5050 2339
rect 4774 2254 4802 2282
rect 5110 2310 5138 2338
rect 5614 2254 5642 2282
rect 6398 2926 6426 2954
rect 7074 4717 7102 4718
rect 7074 4691 7075 4717
rect 7075 4691 7101 4717
rect 7101 4691 7102 4717
rect 7074 4690 7102 4691
rect 7126 4717 7154 4718
rect 7126 4691 7127 4717
rect 7127 4691 7153 4717
rect 7153 4691 7154 4717
rect 7126 4690 7154 4691
rect 7178 4717 7206 4718
rect 7178 4691 7179 4717
rect 7179 4691 7205 4717
rect 7205 4691 7206 4717
rect 7178 4690 7206 4691
rect 6958 4438 6986 4466
rect 6734 4102 6762 4130
rect 6454 2422 6482 2450
rect 6678 2534 6706 2562
rect 6342 2254 6370 2282
rect 5278 2169 5306 2170
rect 5278 2143 5279 2169
rect 5279 2143 5305 2169
rect 5305 2143 5306 2169
rect 5278 2142 5306 2143
rect 6622 2254 6650 2282
rect 6622 2142 6650 2170
rect 5996 1973 6024 1974
rect 5996 1947 5997 1973
rect 5997 1947 6023 1973
rect 6023 1947 6024 1973
rect 5996 1946 6024 1947
rect 6048 1973 6076 1974
rect 6048 1947 6049 1973
rect 6049 1947 6075 1973
rect 6075 1947 6076 1973
rect 6048 1946 6076 1947
rect 6100 1973 6128 1974
rect 6100 1947 6101 1973
rect 6101 1947 6127 1973
rect 6127 1947 6128 1973
rect 6100 1946 6128 1947
rect 6958 3374 6986 3402
rect 6846 2534 6874 2562
rect 7074 3933 7102 3934
rect 7074 3907 7075 3933
rect 7075 3907 7101 3933
rect 7101 3907 7102 3933
rect 7074 3906 7102 3907
rect 7126 3933 7154 3934
rect 7126 3907 7127 3933
rect 7127 3907 7153 3933
rect 7153 3907 7154 3933
rect 7126 3906 7154 3907
rect 7178 3933 7206 3934
rect 7178 3907 7179 3933
rect 7179 3907 7205 3933
rect 7205 3907 7206 3933
rect 7178 3906 7206 3907
rect 7350 3822 7378 3850
rect 7014 3486 7042 3514
rect 6958 2953 6986 2954
rect 6958 2927 6959 2953
rect 6959 2927 6985 2953
rect 6985 2927 6986 2953
rect 6958 2926 6986 2927
rect 6958 2758 6986 2786
rect 7070 3766 7098 3794
rect 7074 3149 7102 3150
rect 7074 3123 7075 3149
rect 7075 3123 7101 3149
rect 7101 3123 7102 3149
rect 7074 3122 7102 3123
rect 7126 3149 7154 3150
rect 7126 3123 7127 3149
rect 7127 3123 7153 3149
rect 7153 3123 7154 3149
rect 7126 3122 7154 3123
rect 7178 3149 7206 3150
rect 7178 3123 7179 3149
rect 7179 3123 7205 3149
rect 7205 3123 7206 3149
rect 7178 3122 7206 3123
rect 7294 3486 7322 3514
rect 7854 5614 7882 5642
rect 7910 5558 7938 5586
rect 8022 6006 8050 6034
rect 8152 5893 8180 5894
rect 8152 5867 8153 5893
rect 8153 5867 8179 5893
rect 8179 5867 8180 5893
rect 8152 5866 8180 5867
rect 8204 5893 8232 5894
rect 8204 5867 8205 5893
rect 8205 5867 8231 5893
rect 8231 5867 8232 5893
rect 8204 5866 8232 5867
rect 8256 5893 8284 5894
rect 8256 5867 8257 5893
rect 8257 5867 8283 5893
rect 8283 5867 8284 5893
rect 8256 5866 8284 5867
rect 8750 6033 8778 6034
rect 8750 6007 8751 6033
rect 8751 6007 8777 6033
rect 8777 6007 8778 6033
rect 8750 6006 8778 6007
rect 8358 5782 8386 5810
rect 8750 5782 8778 5810
rect 9086 7630 9114 7658
rect 8862 6873 8890 6874
rect 8862 6847 8863 6873
rect 8863 6847 8889 6873
rect 8889 6847 8890 6873
rect 8862 6846 8890 6847
rect 8806 5726 8834 5754
rect 8190 5361 8218 5362
rect 8190 5335 8191 5361
rect 8191 5335 8217 5361
rect 8217 5335 8218 5361
rect 8190 5334 8218 5335
rect 8134 5305 8162 5306
rect 8134 5279 8135 5305
rect 8135 5279 8161 5305
rect 8161 5279 8162 5305
rect 8134 5278 8162 5279
rect 7910 4857 7938 4858
rect 7910 4831 7911 4857
rect 7911 4831 7937 4857
rect 7937 4831 7938 4857
rect 7910 4830 7938 4831
rect 7462 3766 7490 3794
rect 7462 3430 7490 3458
rect 7518 3318 7546 3346
rect 7406 2982 7434 3010
rect 7238 2758 7266 2786
rect 7910 4158 7938 4186
rect 8152 5109 8180 5110
rect 8152 5083 8153 5109
rect 8153 5083 8179 5109
rect 8179 5083 8180 5109
rect 8152 5082 8180 5083
rect 8204 5109 8232 5110
rect 8204 5083 8205 5109
rect 8205 5083 8231 5109
rect 8231 5083 8232 5109
rect 8204 5082 8232 5083
rect 8256 5109 8284 5110
rect 8256 5083 8257 5109
rect 8257 5083 8283 5109
rect 8283 5083 8284 5109
rect 8256 5082 8284 5083
rect 8302 4998 8330 5026
rect 8358 4550 8386 4578
rect 8358 4438 8386 4466
rect 8152 4325 8180 4326
rect 8152 4299 8153 4325
rect 8153 4299 8179 4325
rect 8179 4299 8180 4325
rect 8152 4298 8180 4299
rect 8204 4325 8232 4326
rect 8204 4299 8205 4325
rect 8205 4299 8231 4325
rect 8231 4299 8232 4325
rect 8204 4298 8232 4299
rect 8256 4325 8284 4326
rect 8256 4299 8257 4325
rect 8257 4299 8283 4325
rect 8283 4299 8284 4325
rect 8256 4298 8284 4299
rect 9086 5782 9114 5810
rect 9230 7069 9258 7070
rect 9230 7043 9231 7069
rect 9231 7043 9257 7069
rect 9257 7043 9258 7069
rect 9230 7042 9258 7043
rect 9282 7069 9310 7070
rect 9282 7043 9283 7069
rect 9283 7043 9309 7069
rect 9309 7043 9310 7069
rect 9282 7042 9310 7043
rect 9334 7069 9362 7070
rect 9334 7043 9335 7069
rect 9335 7043 9361 7069
rect 9361 7043 9362 7069
rect 9334 7042 9362 7043
rect 9230 6285 9258 6286
rect 9230 6259 9231 6285
rect 9231 6259 9257 6285
rect 9257 6259 9258 6285
rect 9230 6258 9258 6259
rect 9282 6285 9310 6286
rect 9282 6259 9283 6285
rect 9283 6259 9309 6285
rect 9309 6259 9310 6285
rect 9282 6258 9310 6259
rect 9334 6285 9362 6286
rect 9334 6259 9335 6285
rect 9335 6259 9361 6285
rect 9361 6259 9362 6285
rect 9334 6258 9362 6259
rect 8918 5054 8946 5082
rect 9230 5501 9258 5502
rect 9230 5475 9231 5501
rect 9231 5475 9257 5501
rect 9257 5475 9258 5501
rect 9230 5474 9258 5475
rect 9282 5501 9310 5502
rect 9282 5475 9283 5501
rect 9283 5475 9309 5501
rect 9309 5475 9310 5501
rect 9282 5474 9310 5475
rect 9334 5501 9362 5502
rect 9334 5475 9335 5501
rect 9335 5475 9361 5501
rect 9361 5475 9362 5501
rect 9334 5474 9362 5475
rect 8750 4830 8778 4858
rect 8694 4577 8722 4578
rect 8694 4551 8695 4577
rect 8695 4551 8721 4577
rect 8721 4551 8722 4577
rect 8694 4550 8722 4551
rect 9230 4717 9258 4718
rect 9230 4691 9231 4717
rect 9231 4691 9257 4717
rect 9257 4691 9258 4717
rect 9230 4690 9258 4691
rect 9282 4717 9310 4718
rect 9282 4691 9283 4717
rect 9283 4691 9309 4717
rect 9309 4691 9310 4717
rect 9282 4690 9310 4691
rect 9334 4717 9362 4718
rect 9334 4691 9335 4717
rect 9335 4691 9361 4717
rect 9361 4691 9362 4717
rect 9334 4690 9362 4691
rect 8918 3822 8946 3850
rect 8694 3766 8722 3794
rect 8246 3737 8274 3738
rect 8246 3711 8247 3737
rect 8247 3711 8273 3737
rect 8273 3711 8274 3737
rect 8246 3710 8274 3711
rect 8358 3598 8386 3626
rect 8152 3541 8180 3542
rect 8152 3515 8153 3541
rect 8153 3515 8179 3541
rect 8179 3515 8180 3541
rect 8152 3514 8180 3515
rect 8204 3541 8232 3542
rect 8204 3515 8205 3541
rect 8205 3515 8231 3541
rect 8231 3515 8232 3541
rect 8204 3514 8232 3515
rect 8256 3541 8284 3542
rect 8256 3515 8257 3541
rect 8257 3515 8283 3541
rect 8283 3515 8284 3541
rect 8256 3514 8284 3515
rect 8022 3345 8050 3346
rect 8022 3319 8023 3345
rect 8023 3319 8049 3345
rect 8049 3319 8050 3345
rect 8022 3318 8050 3319
rect 8078 3038 8106 3066
rect 7686 2926 7714 2954
rect 7126 2590 7154 2618
rect 7686 2534 7714 2562
rect 6846 2449 6874 2450
rect 6846 2423 6847 2449
rect 6847 2423 6873 2449
rect 6873 2423 6874 2449
rect 6846 2422 6874 2423
rect 6734 2310 6762 2338
rect 7238 2478 7266 2506
rect 6678 2086 6706 2114
rect 6174 1833 6202 1834
rect 6174 1807 6175 1833
rect 6175 1807 6201 1833
rect 6201 1807 6202 1833
rect 6174 1806 6202 1807
rect 4102 1750 4130 1778
rect 5054 1777 5082 1778
rect 5054 1751 5055 1777
rect 5055 1751 5081 1777
rect 5081 1751 5082 1777
rect 5054 1750 5082 1751
rect 6622 1750 6650 1778
rect 7074 2365 7102 2366
rect 7074 2339 7075 2365
rect 7075 2339 7101 2365
rect 7101 2339 7102 2365
rect 7074 2338 7102 2339
rect 7126 2365 7154 2366
rect 7126 2339 7127 2365
rect 7127 2339 7153 2365
rect 7153 2339 7154 2365
rect 7126 2338 7154 2339
rect 7178 2365 7206 2366
rect 7178 2339 7179 2365
rect 7179 2339 7205 2365
rect 7205 2339 7206 2365
rect 7178 2338 7206 2339
rect 8638 3430 8666 3458
rect 8152 2757 8180 2758
rect 8152 2731 8153 2757
rect 8153 2731 8179 2757
rect 8179 2731 8180 2757
rect 8152 2730 8180 2731
rect 8204 2757 8232 2758
rect 8204 2731 8205 2757
rect 8205 2731 8231 2757
rect 8231 2731 8232 2757
rect 8204 2730 8232 2731
rect 8256 2757 8284 2758
rect 8256 2731 8257 2757
rect 8257 2731 8283 2757
rect 8283 2731 8284 2757
rect 8256 2730 8284 2731
rect 8806 2561 8834 2562
rect 8806 2535 8807 2561
rect 8807 2535 8833 2561
rect 8833 2535 8834 2561
rect 8806 2534 8834 2535
rect 8974 3793 9002 3794
rect 8974 3767 8975 3793
rect 8975 3767 9001 3793
rect 9001 3767 9002 3793
rect 8974 3766 9002 3767
rect 9230 3933 9258 3934
rect 9230 3907 9231 3933
rect 9231 3907 9257 3933
rect 9257 3907 9258 3933
rect 9230 3906 9258 3907
rect 9282 3933 9310 3934
rect 9282 3907 9283 3933
rect 9283 3907 9309 3933
rect 9309 3907 9310 3933
rect 9282 3906 9310 3907
rect 9334 3933 9362 3934
rect 9334 3907 9335 3933
rect 9335 3907 9361 3933
rect 9361 3907 9362 3933
rect 9334 3906 9362 3907
rect 9142 3737 9170 3738
rect 9142 3711 9143 3737
rect 9143 3711 9169 3737
rect 9169 3711 9170 3737
rect 9142 3710 9170 3711
rect 9030 3598 9058 3626
rect 9230 3149 9258 3150
rect 9230 3123 9231 3149
rect 9231 3123 9257 3149
rect 9257 3123 9258 3149
rect 9230 3122 9258 3123
rect 9282 3149 9310 3150
rect 9282 3123 9283 3149
rect 9283 3123 9309 3149
rect 9309 3123 9310 3149
rect 9282 3122 9310 3123
rect 9334 3149 9362 3150
rect 9334 3123 9335 3149
rect 9335 3123 9361 3149
rect 9361 3123 9362 3149
rect 9334 3122 9362 3123
rect 9142 2590 9170 2618
rect 9230 2365 9258 2366
rect 9230 2339 9231 2365
rect 9231 2339 9257 2365
rect 9257 2339 9258 2365
rect 9230 2338 9258 2339
rect 9282 2365 9310 2366
rect 9282 2339 9283 2365
rect 9283 2339 9309 2365
rect 9309 2339 9310 2365
rect 9282 2338 9310 2339
rect 9334 2365 9362 2366
rect 9334 2339 9335 2365
rect 9335 2339 9361 2365
rect 9361 2339 9362 2365
rect 9334 2338 9362 2339
rect 8862 2254 8890 2282
rect 8694 2113 8722 2114
rect 8694 2087 8695 2113
rect 8695 2087 8721 2113
rect 8721 2087 8722 2113
rect 8694 2086 8722 2087
rect 8152 1973 8180 1974
rect 8152 1947 8153 1973
rect 8153 1947 8179 1973
rect 8179 1947 8180 1973
rect 8152 1946 8180 1947
rect 8204 1973 8232 1974
rect 8204 1947 8205 1973
rect 8205 1947 8231 1973
rect 8231 1947 8232 1973
rect 8204 1946 8232 1947
rect 8256 1973 8284 1974
rect 8256 1947 8257 1973
rect 8257 1947 8283 1973
rect 8283 1947 8284 1973
rect 8256 1946 8284 1947
rect 7350 1750 7378 1778
rect 2762 1581 2790 1582
rect 2762 1555 2763 1581
rect 2763 1555 2789 1581
rect 2789 1555 2790 1581
rect 2762 1554 2790 1555
rect 2814 1581 2842 1582
rect 2814 1555 2815 1581
rect 2815 1555 2841 1581
rect 2841 1555 2842 1581
rect 2814 1554 2842 1555
rect 2866 1581 2894 1582
rect 2866 1555 2867 1581
rect 2867 1555 2893 1581
rect 2893 1555 2894 1581
rect 2866 1554 2894 1555
rect 4918 1581 4946 1582
rect 4918 1555 4919 1581
rect 4919 1555 4945 1581
rect 4945 1555 4946 1581
rect 4918 1554 4946 1555
rect 4970 1581 4998 1582
rect 4970 1555 4971 1581
rect 4971 1555 4997 1581
rect 4997 1555 4998 1581
rect 4970 1554 4998 1555
rect 5022 1581 5050 1582
rect 5022 1555 5023 1581
rect 5023 1555 5049 1581
rect 5049 1555 5050 1581
rect 5022 1554 5050 1555
rect 7074 1581 7102 1582
rect 7074 1555 7075 1581
rect 7075 1555 7101 1581
rect 7101 1555 7102 1581
rect 7074 1554 7102 1555
rect 7126 1581 7154 1582
rect 7126 1555 7127 1581
rect 7127 1555 7153 1581
rect 7153 1555 7154 1581
rect 7126 1554 7154 1555
rect 7178 1581 7206 1582
rect 7178 1555 7179 1581
rect 7179 1555 7205 1581
rect 7205 1555 7206 1581
rect 7178 1554 7206 1555
rect 966 1246 994 1274
rect 9230 1581 9258 1582
rect 9230 1555 9231 1581
rect 9231 1555 9257 1581
rect 9257 1555 9258 1581
rect 9230 1554 9258 1555
rect 9282 1581 9310 1582
rect 9282 1555 9283 1581
rect 9283 1555 9309 1581
rect 9309 1555 9310 1581
rect 9282 1554 9310 1555
rect 9334 1581 9362 1582
rect 9334 1555 9335 1581
rect 9335 1555 9361 1581
rect 9361 1555 9362 1581
rect 9334 1554 9362 1555
rect 9086 574 9114 602
<< metal3 >>
rect 9600 9226 10000 9240
rect 7905 9198 7910 9226
rect 7938 9198 10000 9226
rect 9600 9184 10000 9198
rect 0 8666 400 8680
rect 0 8638 854 8666
rect 882 8638 887 8666
rect 0 8624 400 8638
rect 7401 8358 7406 8386
rect 7434 8358 8582 8386
rect 8610 8358 8615 8386
rect 1679 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1821 8246
rect 3835 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3977 8246
rect 5991 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6133 8246
rect 8147 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8289 8246
rect 849 8078 854 8106
rect 882 8078 1246 8106
rect 1274 8078 1279 8106
rect 8577 8078 8582 8106
rect 8610 8078 8862 8106
rect 8890 8078 8895 8106
rect 8185 8022 8190 8050
rect 8218 8022 8806 8050
rect 8834 8022 8839 8050
rect 9600 7994 10000 8008
rect 5441 7966 5446 7994
rect 5474 7966 6118 7994
rect 6146 7966 6151 7994
rect 7401 7966 7406 7994
rect 7434 7966 10000 7994
rect 9600 7952 10000 7966
rect 1017 7910 1022 7938
rect 1050 7910 1862 7938
rect 1890 7910 1895 7938
rect 2757 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2899 7854
rect 4913 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5055 7854
rect 7069 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7211 7854
rect 9225 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9367 7854
rect 3425 7630 3430 7658
rect 3458 7630 5782 7658
rect 5810 7630 5815 7658
rect 6897 7630 6902 7658
rect 6930 7630 7574 7658
rect 7602 7630 7607 7658
rect 8409 7630 8414 7658
rect 8442 7630 9086 7658
rect 9114 7630 9119 7658
rect 4937 7574 4942 7602
rect 4970 7574 5446 7602
rect 5474 7574 5479 7602
rect 6225 7574 6230 7602
rect 6258 7574 6510 7602
rect 6538 7574 6543 7602
rect 4489 7462 4494 7490
rect 4522 7462 4774 7490
rect 4802 7462 4998 7490
rect 5026 7462 5031 7490
rect 1679 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1821 7462
rect 3835 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3977 7462
rect 5991 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6133 7462
rect 8147 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8289 7462
rect 3089 7350 3094 7378
rect 3122 7350 3598 7378
rect 3626 7350 4326 7378
rect 4354 7350 4359 7378
rect 5273 7238 5278 7266
rect 5306 7238 5894 7266
rect 5922 7238 6398 7266
rect 6426 7238 6431 7266
rect 7233 7238 7238 7266
rect 7266 7238 8750 7266
rect 8778 7238 8783 7266
rect 4657 7182 4662 7210
rect 4690 7182 5558 7210
rect 5586 7182 5591 7210
rect 6449 7182 6454 7210
rect 6482 7182 7126 7210
rect 7154 7182 7159 7210
rect 7513 7182 7518 7210
rect 7546 7182 7966 7210
rect 7994 7182 7999 7210
rect 3369 7126 3374 7154
rect 3402 7126 3934 7154
rect 3962 7126 4774 7154
rect 4802 7126 4807 7154
rect 5161 7126 5166 7154
rect 5194 7126 5199 7154
rect 5665 7126 5670 7154
rect 5698 7126 5838 7154
rect 5866 7126 5871 7154
rect 6001 7126 6006 7154
rect 6034 7126 6678 7154
rect 6706 7126 6711 7154
rect 2757 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2899 7070
rect 4774 6986 4802 7126
rect 4913 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5055 7070
rect 5166 7042 5194 7126
rect 7069 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7211 7070
rect 9225 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9367 7070
rect 5166 7014 5894 7042
rect 5922 7014 5927 7042
rect 4774 6958 4998 6986
rect 5026 6958 5031 6986
rect 5833 6958 5838 6986
rect 5866 6958 5871 6986
rect 4489 6902 4494 6930
rect 4522 6902 5166 6930
rect 5194 6902 5199 6930
rect 5838 6874 5866 6958
rect 5838 6846 5950 6874
rect 5978 6846 5983 6874
rect 6169 6846 6174 6874
rect 6202 6846 6510 6874
rect 6538 6846 6543 6874
rect 8409 6846 8414 6874
rect 8442 6846 8862 6874
rect 8890 6846 8895 6874
rect 2977 6790 2982 6818
rect 3010 6790 5222 6818
rect 5250 6790 5255 6818
rect 9600 6762 10000 6776
rect 4041 6734 4046 6762
rect 4074 6734 4438 6762
rect 4466 6734 4718 6762
rect 4746 6734 5110 6762
rect 5138 6734 5143 6762
rect 5894 6734 6062 6762
rect 6090 6734 6986 6762
rect 7905 6734 7910 6762
rect 7938 6734 10000 6762
rect 5894 6706 5922 6734
rect 5777 6678 5782 6706
rect 5810 6678 5922 6706
rect 1679 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1821 6678
rect 3835 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3977 6678
rect 5991 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6133 6678
rect 6958 6650 6986 6734
rect 9600 6720 10000 6734
rect 8147 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8289 6678
rect 5329 6622 5334 6650
rect 5362 6622 5390 6650
rect 5418 6622 5423 6650
rect 6953 6622 6958 6650
rect 6986 6622 7294 6650
rect 7322 6622 7327 6650
rect 4657 6566 4662 6594
rect 4690 6566 5278 6594
rect 5306 6566 5311 6594
rect 6169 6566 6174 6594
rect 6202 6566 6566 6594
rect 6594 6566 6599 6594
rect 4377 6510 4382 6538
rect 4410 6510 4415 6538
rect 4601 6510 4606 6538
rect 4634 6510 5334 6538
rect 5362 6510 5502 6538
rect 5530 6510 5535 6538
rect 7401 6510 7406 6538
rect 7434 6510 8022 6538
rect 8050 6510 8055 6538
rect 4382 6482 4410 6510
rect 4209 6454 4214 6482
rect 4242 6454 5306 6482
rect 5889 6454 5894 6482
rect 5922 6454 6006 6482
rect 6034 6454 6039 6482
rect 7009 6454 7014 6482
rect 7042 6454 8470 6482
rect 8498 6454 8503 6482
rect 5278 6426 5306 6454
rect 4041 6398 4046 6426
rect 4074 6398 4270 6426
rect 4298 6398 4606 6426
rect 4634 6398 4639 6426
rect 5273 6398 5278 6426
rect 5306 6398 6174 6426
rect 6202 6398 6207 6426
rect 7289 6398 7294 6426
rect 7322 6398 8694 6426
rect 8722 6398 8727 6426
rect 5278 6342 5670 6370
rect 5698 6342 5703 6370
rect 6953 6342 6958 6370
rect 6986 6342 7126 6370
rect 7154 6342 7378 6370
rect 5278 6314 5306 6342
rect 5273 6286 5278 6314
rect 5306 6286 5311 6314
rect 5553 6286 5558 6314
rect 5586 6286 6062 6314
rect 6090 6286 6095 6314
rect 2757 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2899 6286
rect 4913 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5055 6286
rect 7069 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7211 6286
rect 7350 6258 7378 6342
rect 9225 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9367 6286
rect 5161 6230 5166 6258
rect 5194 6230 5838 6258
rect 5866 6230 5871 6258
rect 7345 6230 7350 6258
rect 7378 6230 7383 6258
rect 0 6202 400 6216
rect 0 6174 854 6202
rect 882 6174 1246 6202
rect 1274 6174 1279 6202
rect 2473 6174 2478 6202
rect 2506 6174 4830 6202
rect 4858 6174 5054 6202
rect 5082 6174 5087 6202
rect 5371 6174 5390 6202
rect 5418 6174 5423 6202
rect 0 6160 400 6174
rect 4321 6118 4326 6146
rect 4354 6118 4662 6146
rect 4690 6118 4695 6146
rect 6897 6118 6902 6146
rect 6930 6118 8638 6146
rect 8666 6118 8671 6146
rect 1969 6062 1974 6090
rect 2002 6062 2702 6090
rect 2730 6062 2735 6090
rect 3985 6062 3990 6090
rect 4018 6062 4382 6090
rect 4410 6062 4415 6090
rect 5945 6062 5950 6090
rect 5978 6062 6566 6090
rect 6594 6062 7966 6090
rect 7994 6062 7999 6090
rect 5721 6006 5726 6034
rect 5754 6006 6062 6034
rect 6090 6006 6095 6034
rect 8017 6006 8022 6034
rect 8050 6006 8750 6034
rect 8778 6006 8783 6034
rect 2305 5950 2310 5978
rect 2338 5950 4942 5978
rect 4970 5950 4975 5978
rect 5273 5950 5278 5978
rect 5306 5950 5894 5978
rect 5922 5950 5927 5978
rect 6001 5950 6006 5978
rect 6034 5950 6202 5978
rect 1679 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1821 5894
rect 3835 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3977 5894
rect 5991 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6133 5894
rect 6174 5866 6202 5950
rect 8147 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8289 5894
rect 6174 5838 7182 5866
rect 7210 5838 7215 5866
rect 5161 5782 5166 5810
rect 5194 5782 6286 5810
rect 6314 5782 6319 5810
rect 8353 5782 8358 5810
rect 8386 5782 8750 5810
rect 8778 5782 9086 5810
rect 9114 5782 9119 5810
rect 7289 5726 7294 5754
rect 7322 5726 8806 5754
rect 8834 5726 8839 5754
rect 4545 5670 4550 5698
rect 4578 5670 4886 5698
rect 4914 5670 4919 5698
rect 4993 5670 4998 5698
rect 5026 5670 5110 5698
rect 5138 5670 5950 5698
rect 5978 5670 5983 5698
rect 5166 5614 6734 5642
rect 6762 5614 6767 5642
rect 7065 5614 7070 5642
rect 7098 5614 7406 5642
rect 7434 5614 7854 5642
rect 7882 5614 7887 5642
rect 5166 5586 5194 5614
rect 6342 5586 6370 5614
rect 1638 5558 5166 5586
rect 5194 5558 5199 5586
rect 5665 5558 5670 5586
rect 5698 5558 6174 5586
rect 6202 5558 6207 5586
rect 6337 5558 6342 5586
rect 6370 5558 6375 5586
rect 7905 5558 7910 5586
rect 7938 5558 9450 5586
rect 1638 5474 1666 5558
rect 9422 5530 9450 5558
rect 9600 5530 10000 5544
rect 5945 5502 5950 5530
rect 5978 5502 6230 5530
rect 6258 5502 6263 5530
rect 9422 5502 10000 5530
rect 2757 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2899 5502
rect 4913 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5055 5502
rect 7069 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7211 5502
rect 9225 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9367 5502
rect 9600 5488 10000 5502
rect 1633 5446 1638 5474
rect 1666 5446 1671 5474
rect 5329 5446 5334 5474
rect 5362 5446 6930 5474
rect 6902 5418 6930 5446
rect 3313 5390 3318 5418
rect 3346 5390 6734 5418
rect 6762 5390 6767 5418
rect 6902 5390 7182 5418
rect 7210 5390 7215 5418
rect 4433 5334 4438 5362
rect 4466 5334 4774 5362
rect 4802 5334 4807 5362
rect 5329 5334 5334 5362
rect 5362 5334 5614 5362
rect 5642 5334 8190 5362
rect 8218 5334 8223 5362
rect 2585 5278 2590 5306
rect 2618 5278 3486 5306
rect 3514 5278 3519 5306
rect 3593 5278 3598 5306
rect 3626 5278 4550 5306
rect 4578 5278 4830 5306
rect 4858 5278 4863 5306
rect 4937 5278 4942 5306
rect 4970 5278 5222 5306
rect 5250 5278 5255 5306
rect 7457 5278 7462 5306
rect 7490 5278 8134 5306
rect 8162 5278 8167 5306
rect 2865 5222 2870 5250
rect 2898 5222 3710 5250
rect 3738 5222 3743 5250
rect 3929 5222 3934 5250
rect 3962 5222 4102 5250
rect 4130 5222 4135 5250
rect 4265 5222 4270 5250
rect 4298 5222 5446 5250
rect 5474 5222 5479 5250
rect 4041 5166 4046 5194
rect 4074 5166 4774 5194
rect 4802 5166 4807 5194
rect 1679 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1821 5110
rect 3835 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3977 5110
rect 5991 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6133 5110
rect 8147 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8289 5110
rect 3089 5054 3094 5082
rect 3122 5054 3318 5082
rect 3346 5054 3351 5082
rect 4097 5054 4102 5082
rect 4130 5054 5642 5082
rect 2697 4998 2702 5026
rect 2730 4998 2982 5026
rect 3010 4998 3015 5026
rect 5614 4970 5642 5054
rect 8358 5054 8918 5082
rect 8946 5054 8951 5082
rect 8358 5026 8386 5054
rect 5721 4998 5726 5026
rect 5754 4998 6174 5026
rect 6202 4998 6207 5026
rect 8297 4998 8302 5026
rect 8330 4998 8386 5026
rect 3033 4942 3038 4970
rect 3066 4942 3654 4970
rect 3682 4942 4550 4970
rect 4578 4942 4583 4970
rect 5614 4942 6118 4970
rect 6146 4942 6151 4970
rect 7905 4830 7910 4858
rect 7938 4830 8750 4858
rect 8778 4830 8783 4858
rect 2757 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2899 4718
rect 4913 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5055 4718
rect 7069 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7211 4718
rect 9225 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9367 4718
rect 3201 4606 3206 4634
rect 3234 4606 3710 4634
rect 3738 4606 3743 4634
rect 2137 4550 2142 4578
rect 2170 4550 2534 4578
rect 2562 4550 2758 4578
rect 2786 4550 2791 4578
rect 8353 4550 8358 4578
rect 8386 4550 8694 4578
rect 8722 4550 8727 4578
rect 2865 4494 2870 4522
rect 2898 4494 3038 4522
rect 3066 4494 3071 4522
rect 5385 4438 5390 4466
rect 5418 4438 5894 4466
rect 5922 4438 5927 4466
rect 6953 4438 6958 4466
rect 6986 4438 8358 4466
rect 8386 4438 8391 4466
rect 1679 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1821 4326
rect 3835 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3977 4326
rect 5991 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6133 4326
rect 8147 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8289 4326
rect 9600 4298 10000 4312
rect 8358 4270 10000 4298
rect 8358 4186 8386 4270
rect 9600 4256 10000 4270
rect 7905 4158 7910 4186
rect 7938 4158 8386 4186
rect 6001 4102 6006 4130
rect 6034 4102 6286 4130
rect 6314 4102 6734 4130
rect 6762 4102 6767 4130
rect 1745 4046 1750 4074
rect 1778 4046 1862 4074
rect 1890 4046 1895 4074
rect 4489 4046 4494 4074
rect 4522 4046 4942 4074
rect 4970 4046 5502 4074
rect 5530 4046 5535 4074
rect 3873 3990 3878 4018
rect 3906 3990 4438 4018
rect 4466 3990 5222 4018
rect 5250 3990 5894 4018
rect 5922 3990 5927 4018
rect 2757 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2899 3934
rect 4913 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5055 3934
rect 7069 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7211 3934
rect 9225 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9367 3934
rect 2963 3822 2982 3850
rect 3010 3822 7350 3850
rect 7378 3822 8918 3850
rect 8946 3822 8951 3850
rect 1017 3766 1022 3794
rect 1050 3766 1302 3794
rect 1330 3766 1862 3794
rect 1890 3766 1895 3794
rect 2473 3766 2478 3794
rect 2506 3766 3094 3794
rect 3122 3766 3127 3794
rect 7065 3766 7070 3794
rect 7098 3766 7462 3794
rect 7490 3766 7495 3794
rect 8689 3766 8694 3794
rect 8722 3766 8974 3794
rect 9002 3766 9007 3794
rect 0 3738 400 3752
rect 0 3710 910 3738
rect 938 3710 943 3738
rect 1073 3710 1078 3738
rect 1106 3710 2310 3738
rect 2338 3710 2343 3738
rect 3145 3710 3150 3738
rect 3178 3710 3654 3738
rect 3682 3710 3822 3738
rect 3850 3710 3855 3738
rect 8241 3710 8246 3738
rect 8274 3710 9142 3738
rect 9170 3710 9175 3738
rect 0 3696 400 3710
rect 1409 3654 1414 3682
rect 1442 3654 1750 3682
rect 1778 3654 2198 3682
rect 2226 3654 2231 3682
rect 8353 3598 8358 3626
rect 8386 3598 9030 3626
rect 9058 3598 9063 3626
rect 1679 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1821 3542
rect 3835 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3977 3542
rect 5991 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6133 3542
rect 8147 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8289 3542
rect 2025 3486 2030 3514
rect 2058 3486 2534 3514
rect 2562 3486 3038 3514
rect 3066 3486 3071 3514
rect 7009 3486 7014 3514
rect 7042 3486 7294 3514
rect 7322 3486 7327 3514
rect 2193 3430 2198 3458
rect 2226 3430 3094 3458
rect 3122 3430 3127 3458
rect 7457 3430 7462 3458
rect 7490 3430 8638 3458
rect 8666 3430 8671 3458
rect 1521 3374 1526 3402
rect 1554 3374 2254 3402
rect 2282 3374 2287 3402
rect 5273 3374 5278 3402
rect 5306 3374 6062 3402
rect 6090 3374 6958 3402
rect 6986 3374 6991 3402
rect 3649 3318 3654 3346
rect 3682 3318 3934 3346
rect 3962 3318 3967 3346
rect 7513 3318 7518 3346
rect 7546 3318 8022 3346
rect 8050 3318 8055 3346
rect 1297 3262 1302 3290
rect 1330 3262 1918 3290
rect 1946 3262 1951 3290
rect 4209 3262 4214 3290
rect 4242 3262 4998 3290
rect 5026 3262 5031 3290
rect 2757 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2899 3150
rect 4913 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5055 3150
rect 7069 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7211 3150
rect 9225 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9367 3150
rect 3486 3094 4270 3122
rect 4298 3094 4303 3122
rect 3486 3066 3514 3094
rect 9600 3066 10000 3080
rect 2697 3038 2702 3066
rect 2730 3038 3094 3066
rect 3122 3038 3486 3066
rect 3514 3038 3519 3066
rect 4153 3038 4158 3066
rect 4186 3038 5222 3066
rect 5250 3038 5255 3066
rect 8073 3038 8078 3066
rect 8106 3038 10000 3066
rect 9600 3024 10000 3038
rect 4377 2982 4382 3010
rect 4410 2982 4998 3010
rect 5026 2982 7406 3010
rect 7434 2982 7439 3010
rect 1129 2926 1134 2954
rect 1162 2926 2142 2954
rect 2170 2926 2814 2954
rect 2842 2926 3710 2954
rect 3738 2926 3743 2954
rect 6393 2926 6398 2954
rect 6426 2926 6958 2954
rect 6986 2926 7686 2954
rect 7714 2926 7719 2954
rect 3201 2870 3206 2898
rect 3234 2870 3766 2898
rect 3794 2870 3799 2898
rect 3985 2870 3990 2898
rect 4018 2870 6230 2898
rect 6258 2870 6263 2898
rect 4041 2814 4046 2842
rect 4074 2814 4886 2842
rect 4914 2814 4919 2842
rect 6953 2758 6958 2786
rect 6986 2758 7238 2786
rect 7266 2758 7271 2786
rect 1679 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1821 2758
rect 3835 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3977 2758
rect 5991 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6133 2758
rect 8147 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8289 2758
rect 3313 2646 3318 2674
rect 3346 2646 3878 2674
rect 3906 2646 3911 2674
rect 2473 2590 2478 2618
rect 2506 2590 2926 2618
rect 2954 2590 2959 2618
rect 4993 2590 4998 2618
rect 5026 2590 6006 2618
rect 6034 2590 6039 2618
rect 7121 2590 7126 2618
rect 7154 2590 9142 2618
rect 9170 2590 9175 2618
rect 2585 2534 2590 2562
rect 2618 2534 2982 2562
rect 3010 2534 3015 2562
rect 4321 2534 4326 2562
rect 4354 2534 6678 2562
rect 6706 2534 6711 2562
rect 6841 2534 6846 2562
rect 6874 2534 6879 2562
rect 7681 2534 7686 2562
rect 7714 2534 8806 2562
rect 8834 2534 8839 2562
rect 6846 2506 6874 2534
rect 6846 2478 7238 2506
rect 7266 2478 7271 2506
rect 4713 2422 4718 2450
rect 4746 2422 6454 2450
rect 6482 2422 6846 2450
rect 6874 2422 6879 2450
rect 2757 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2899 2366
rect 4913 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5055 2366
rect 7069 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7211 2366
rect 9225 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9367 2366
rect 5105 2310 5110 2338
rect 5138 2310 6734 2338
rect 6762 2310 6767 2338
rect 4769 2254 4774 2282
rect 4802 2254 5614 2282
rect 5642 2254 6342 2282
rect 6370 2254 6375 2282
rect 6617 2254 6622 2282
rect 6650 2254 8862 2282
rect 8890 2254 8895 2282
rect 3089 2142 3094 2170
rect 3122 2142 3934 2170
rect 3962 2142 3967 2170
rect 5273 2142 5278 2170
rect 5306 2142 6622 2170
rect 6650 2142 6655 2170
rect 6673 2086 6678 2114
rect 6706 2086 8694 2114
rect 8722 2086 8727 2114
rect 1679 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1821 1974
rect 3835 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3977 1974
rect 5991 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6133 1974
rect 8147 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8289 1974
rect 9600 1834 10000 1848
rect 6169 1806 6174 1834
rect 6202 1806 10000 1834
rect 9600 1792 10000 1806
rect 4097 1750 4102 1778
rect 4130 1750 5054 1778
rect 5082 1750 6622 1778
rect 6650 1750 7350 1778
rect 7378 1750 7383 1778
rect 2757 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2899 1582
rect 4913 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5055 1582
rect 7069 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7211 1582
rect 9225 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9367 1582
rect 0 1274 400 1288
rect 0 1246 966 1274
rect 994 1246 999 1274
rect 0 1232 400 1246
rect 9600 602 10000 616
rect 9081 574 9086 602
rect 9114 574 10000 602
rect 9600 560 10000 574
<< via3 >>
rect 1684 8218 1712 8246
rect 1736 8218 1764 8246
rect 1788 8218 1816 8246
rect 3840 8218 3868 8246
rect 3892 8218 3920 8246
rect 3944 8218 3972 8246
rect 5996 8218 6024 8246
rect 6048 8218 6076 8246
rect 6100 8218 6128 8246
rect 8152 8218 8180 8246
rect 8204 8218 8232 8246
rect 8256 8218 8284 8246
rect 2762 7826 2790 7854
rect 2814 7826 2842 7854
rect 2866 7826 2894 7854
rect 4918 7826 4946 7854
rect 4970 7826 4998 7854
rect 5022 7826 5050 7854
rect 7074 7826 7102 7854
rect 7126 7826 7154 7854
rect 7178 7826 7206 7854
rect 9230 7826 9258 7854
rect 9282 7826 9310 7854
rect 9334 7826 9362 7854
rect 1684 7434 1712 7462
rect 1736 7434 1764 7462
rect 1788 7434 1816 7462
rect 3840 7434 3868 7462
rect 3892 7434 3920 7462
rect 3944 7434 3972 7462
rect 5996 7434 6024 7462
rect 6048 7434 6076 7462
rect 6100 7434 6128 7462
rect 8152 7434 8180 7462
rect 8204 7434 8232 7462
rect 8256 7434 8284 7462
rect 2762 7042 2790 7070
rect 2814 7042 2842 7070
rect 2866 7042 2894 7070
rect 4918 7042 4946 7070
rect 4970 7042 4998 7070
rect 5022 7042 5050 7070
rect 7074 7042 7102 7070
rect 7126 7042 7154 7070
rect 7178 7042 7206 7070
rect 9230 7042 9258 7070
rect 9282 7042 9310 7070
rect 9334 7042 9362 7070
rect 5894 7014 5922 7042
rect 1684 6650 1712 6678
rect 1736 6650 1764 6678
rect 1788 6650 1816 6678
rect 3840 6650 3868 6678
rect 3892 6650 3920 6678
rect 3944 6650 3972 6678
rect 5996 6650 6024 6678
rect 6048 6650 6076 6678
rect 6100 6650 6128 6678
rect 8152 6650 8180 6678
rect 8204 6650 8232 6678
rect 8256 6650 8284 6678
rect 5390 6622 5418 6650
rect 5894 6454 5922 6482
rect 2762 6258 2790 6286
rect 2814 6258 2842 6286
rect 2866 6258 2894 6286
rect 4918 6258 4946 6286
rect 4970 6258 4998 6286
rect 5022 6258 5050 6286
rect 7074 6258 7102 6286
rect 7126 6258 7154 6286
rect 7178 6258 7206 6286
rect 9230 6258 9258 6286
rect 9282 6258 9310 6286
rect 9334 6258 9362 6286
rect 5390 6174 5418 6202
rect 1684 5866 1712 5894
rect 1736 5866 1764 5894
rect 1788 5866 1816 5894
rect 3840 5866 3868 5894
rect 3892 5866 3920 5894
rect 3944 5866 3972 5894
rect 5996 5866 6024 5894
rect 6048 5866 6076 5894
rect 6100 5866 6128 5894
rect 8152 5866 8180 5894
rect 8204 5866 8232 5894
rect 8256 5866 8284 5894
rect 2762 5474 2790 5502
rect 2814 5474 2842 5502
rect 2866 5474 2894 5502
rect 4918 5474 4946 5502
rect 4970 5474 4998 5502
rect 5022 5474 5050 5502
rect 7074 5474 7102 5502
rect 7126 5474 7154 5502
rect 7178 5474 7206 5502
rect 9230 5474 9258 5502
rect 9282 5474 9310 5502
rect 9334 5474 9362 5502
rect 1684 5082 1712 5110
rect 1736 5082 1764 5110
rect 1788 5082 1816 5110
rect 3840 5082 3868 5110
rect 3892 5082 3920 5110
rect 3944 5082 3972 5110
rect 5996 5082 6024 5110
rect 6048 5082 6076 5110
rect 6100 5082 6128 5110
rect 8152 5082 8180 5110
rect 8204 5082 8232 5110
rect 8256 5082 8284 5110
rect 2762 4690 2790 4718
rect 2814 4690 2842 4718
rect 2866 4690 2894 4718
rect 4918 4690 4946 4718
rect 4970 4690 4998 4718
rect 5022 4690 5050 4718
rect 7074 4690 7102 4718
rect 7126 4690 7154 4718
rect 7178 4690 7206 4718
rect 9230 4690 9258 4718
rect 9282 4690 9310 4718
rect 9334 4690 9362 4718
rect 1684 4298 1712 4326
rect 1736 4298 1764 4326
rect 1788 4298 1816 4326
rect 3840 4298 3868 4326
rect 3892 4298 3920 4326
rect 3944 4298 3972 4326
rect 5996 4298 6024 4326
rect 6048 4298 6076 4326
rect 6100 4298 6128 4326
rect 8152 4298 8180 4326
rect 8204 4298 8232 4326
rect 8256 4298 8284 4326
rect 2762 3906 2790 3934
rect 2814 3906 2842 3934
rect 2866 3906 2894 3934
rect 4918 3906 4946 3934
rect 4970 3906 4998 3934
rect 5022 3906 5050 3934
rect 7074 3906 7102 3934
rect 7126 3906 7154 3934
rect 7178 3906 7206 3934
rect 9230 3906 9258 3934
rect 9282 3906 9310 3934
rect 9334 3906 9362 3934
rect 2982 3822 3010 3850
rect 1684 3514 1712 3542
rect 1736 3514 1764 3542
rect 1788 3514 1816 3542
rect 3840 3514 3868 3542
rect 3892 3514 3920 3542
rect 3944 3514 3972 3542
rect 5996 3514 6024 3542
rect 6048 3514 6076 3542
rect 6100 3514 6128 3542
rect 8152 3514 8180 3542
rect 8204 3514 8232 3542
rect 8256 3514 8284 3542
rect 2762 3122 2790 3150
rect 2814 3122 2842 3150
rect 2866 3122 2894 3150
rect 4918 3122 4946 3150
rect 4970 3122 4998 3150
rect 5022 3122 5050 3150
rect 7074 3122 7102 3150
rect 7126 3122 7154 3150
rect 7178 3122 7206 3150
rect 9230 3122 9258 3150
rect 9282 3122 9310 3150
rect 9334 3122 9362 3150
rect 1684 2730 1712 2758
rect 1736 2730 1764 2758
rect 1788 2730 1816 2758
rect 3840 2730 3868 2758
rect 3892 2730 3920 2758
rect 3944 2730 3972 2758
rect 5996 2730 6024 2758
rect 6048 2730 6076 2758
rect 6100 2730 6128 2758
rect 8152 2730 8180 2758
rect 8204 2730 8232 2758
rect 8256 2730 8284 2758
rect 2982 2534 3010 2562
rect 2762 2338 2790 2366
rect 2814 2338 2842 2366
rect 2866 2338 2894 2366
rect 4918 2338 4946 2366
rect 4970 2338 4998 2366
rect 5022 2338 5050 2366
rect 7074 2338 7102 2366
rect 7126 2338 7154 2366
rect 7178 2338 7206 2366
rect 9230 2338 9258 2366
rect 9282 2338 9310 2366
rect 9334 2338 9362 2366
rect 1684 1946 1712 1974
rect 1736 1946 1764 1974
rect 1788 1946 1816 1974
rect 3840 1946 3868 1974
rect 3892 1946 3920 1974
rect 3944 1946 3972 1974
rect 5996 1946 6024 1974
rect 6048 1946 6076 1974
rect 6100 1946 6128 1974
rect 8152 1946 8180 1974
rect 8204 1946 8232 1974
rect 8256 1946 8284 1974
rect 2762 1554 2790 1582
rect 2814 1554 2842 1582
rect 2866 1554 2894 1582
rect 4918 1554 4946 1582
rect 4970 1554 4998 1582
rect 5022 1554 5050 1582
rect 7074 1554 7102 1582
rect 7126 1554 7154 1582
rect 7178 1554 7206 1582
rect 9230 1554 9258 1582
rect 9282 1554 9310 1582
rect 9334 1554 9362 1582
<< metal4 >>
rect 1670 8246 1830 8262
rect 1670 8218 1684 8246
rect 1712 8218 1736 8246
rect 1764 8218 1788 8246
rect 1816 8218 1830 8246
rect 1670 7462 1830 8218
rect 1670 7434 1684 7462
rect 1712 7434 1736 7462
rect 1764 7434 1788 7462
rect 1816 7434 1830 7462
rect 1670 6678 1830 7434
rect 1670 6650 1684 6678
rect 1712 6650 1736 6678
rect 1764 6650 1788 6678
rect 1816 6650 1830 6678
rect 1670 5894 1830 6650
rect 1670 5866 1684 5894
rect 1712 5866 1736 5894
rect 1764 5866 1788 5894
rect 1816 5866 1830 5894
rect 1670 5110 1830 5866
rect 1670 5082 1684 5110
rect 1712 5082 1736 5110
rect 1764 5082 1788 5110
rect 1816 5082 1830 5110
rect 1670 4326 1830 5082
rect 1670 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1830 4326
rect 1670 3542 1830 4298
rect 1670 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1830 3542
rect 1670 2758 1830 3514
rect 1670 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1830 2758
rect 1670 1974 1830 2730
rect 1670 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1830 1974
rect 1670 1538 1830 1946
rect 2748 7854 2908 8262
rect 2748 7826 2762 7854
rect 2790 7826 2814 7854
rect 2842 7826 2866 7854
rect 2894 7826 2908 7854
rect 2748 7070 2908 7826
rect 2748 7042 2762 7070
rect 2790 7042 2814 7070
rect 2842 7042 2866 7070
rect 2894 7042 2908 7070
rect 2748 6286 2908 7042
rect 2748 6258 2762 6286
rect 2790 6258 2814 6286
rect 2842 6258 2866 6286
rect 2894 6258 2908 6286
rect 2748 5502 2908 6258
rect 2748 5474 2762 5502
rect 2790 5474 2814 5502
rect 2842 5474 2866 5502
rect 2894 5474 2908 5502
rect 2748 4718 2908 5474
rect 2748 4690 2762 4718
rect 2790 4690 2814 4718
rect 2842 4690 2866 4718
rect 2894 4690 2908 4718
rect 2748 3934 2908 4690
rect 2748 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2908 3934
rect 2748 3150 2908 3906
rect 3826 8246 3986 8262
rect 3826 8218 3840 8246
rect 3868 8218 3892 8246
rect 3920 8218 3944 8246
rect 3972 8218 3986 8246
rect 3826 7462 3986 8218
rect 3826 7434 3840 7462
rect 3868 7434 3892 7462
rect 3920 7434 3944 7462
rect 3972 7434 3986 7462
rect 3826 6678 3986 7434
rect 3826 6650 3840 6678
rect 3868 6650 3892 6678
rect 3920 6650 3944 6678
rect 3972 6650 3986 6678
rect 3826 5894 3986 6650
rect 3826 5866 3840 5894
rect 3868 5866 3892 5894
rect 3920 5866 3944 5894
rect 3972 5866 3986 5894
rect 3826 5110 3986 5866
rect 3826 5082 3840 5110
rect 3868 5082 3892 5110
rect 3920 5082 3944 5110
rect 3972 5082 3986 5110
rect 3826 4326 3986 5082
rect 3826 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3986 4326
rect 2748 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2908 3150
rect 2748 2366 2908 3122
rect 2982 3850 3010 3855
rect 2982 2562 3010 3822
rect 2982 2529 3010 2534
rect 3826 3542 3986 4298
rect 3826 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3986 3542
rect 3826 2758 3986 3514
rect 3826 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3986 2758
rect 2748 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2908 2366
rect 2748 1582 2908 2338
rect 2748 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2908 1582
rect 2748 1538 2908 1554
rect 3826 1974 3986 2730
rect 3826 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3986 1974
rect 3826 1538 3986 1946
rect 4904 7854 5064 8262
rect 4904 7826 4918 7854
rect 4946 7826 4970 7854
rect 4998 7826 5022 7854
rect 5050 7826 5064 7854
rect 4904 7070 5064 7826
rect 4904 7042 4918 7070
rect 4946 7042 4970 7070
rect 4998 7042 5022 7070
rect 5050 7042 5064 7070
rect 5982 8246 6142 8262
rect 5982 8218 5996 8246
rect 6024 8218 6048 8246
rect 6076 8218 6100 8246
rect 6128 8218 6142 8246
rect 5982 7462 6142 8218
rect 5982 7434 5996 7462
rect 6024 7434 6048 7462
rect 6076 7434 6100 7462
rect 6128 7434 6142 7462
rect 4904 6286 5064 7042
rect 5894 7042 5922 7047
rect 4904 6258 4918 6286
rect 4946 6258 4970 6286
rect 4998 6258 5022 6286
rect 5050 6258 5064 6286
rect 4904 5502 5064 6258
rect 5390 6650 5418 6655
rect 5390 6202 5418 6622
rect 5894 6482 5922 7014
rect 5894 6449 5922 6454
rect 5982 6678 6142 7434
rect 5982 6650 5996 6678
rect 6024 6650 6048 6678
rect 6076 6650 6100 6678
rect 6128 6650 6142 6678
rect 5390 6169 5418 6174
rect 4904 5474 4918 5502
rect 4946 5474 4970 5502
rect 4998 5474 5022 5502
rect 5050 5474 5064 5502
rect 4904 4718 5064 5474
rect 4904 4690 4918 4718
rect 4946 4690 4970 4718
rect 4998 4690 5022 4718
rect 5050 4690 5064 4718
rect 4904 3934 5064 4690
rect 4904 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5064 3934
rect 4904 3150 5064 3906
rect 4904 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5064 3150
rect 4904 2366 5064 3122
rect 4904 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5064 2366
rect 4904 1582 5064 2338
rect 4904 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5064 1582
rect 4904 1538 5064 1554
rect 5982 5894 6142 6650
rect 5982 5866 5996 5894
rect 6024 5866 6048 5894
rect 6076 5866 6100 5894
rect 6128 5866 6142 5894
rect 5982 5110 6142 5866
rect 5982 5082 5996 5110
rect 6024 5082 6048 5110
rect 6076 5082 6100 5110
rect 6128 5082 6142 5110
rect 5982 4326 6142 5082
rect 5982 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6142 4326
rect 5982 3542 6142 4298
rect 5982 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6142 3542
rect 5982 2758 6142 3514
rect 5982 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6142 2758
rect 5982 1974 6142 2730
rect 5982 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6142 1974
rect 5982 1538 6142 1946
rect 7060 7854 7220 8262
rect 7060 7826 7074 7854
rect 7102 7826 7126 7854
rect 7154 7826 7178 7854
rect 7206 7826 7220 7854
rect 7060 7070 7220 7826
rect 7060 7042 7074 7070
rect 7102 7042 7126 7070
rect 7154 7042 7178 7070
rect 7206 7042 7220 7070
rect 7060 6286 7220 7042
rect 7060 6258 7074 6286
rect 7102 6258 7126 6286
rect 7154 6258 7178 6286
rect 7206 6258 7220 6286
rect 7060 5502 7220 6258
rect 7060 5474 7074 5502
rect 7102 5474 7126 5502
rect 7154 5474 7178 5502
rect 7206 5474 7220 5502
rect 7060 4718 7220 5474
rect 7060 4690 7074 4718
rect 7102 4690 7126 4718
rect 7154 4690 7178 4718
rect 7206 4690 7220 4718
rect 7060 3934 7220 4690
rect 7060 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7220 3934
rect 7060 3150 7220 3906
rect 7060 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7220 3150
rect 7060 2366 7220 3122
rect 7060 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7220 2366
rect 7060 1582 7220 2338
rect 7060 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7220 1582
rect 7060 1538 7220 1554
rect 8138 8246 8298 8262
rect 8138 8218 8152 8246
rect 8180 8218 8204 8246
rect 8232 8218 8256 8246
rect 8284 8218 8298 8246
rect 8138 7462 8298 8218
rect 8138 7434 8152 7462
rect 8180 7434 8204 7462
rect 8232 7434 8256 7462
rect 8284 7434 8298 7462
rect 8138 6678 8298 7434
rect 8138 6650 8152 6678
rect 8180 6650 8204 6678
rect 8232 6650 8256 6678
rect 8284 6650 8298 6678
rect 8138 5894 8298 6650
rect 8138 5866 8152 5894
rect 8180 5866 8204 5894
rect 8232 5866 8256 5894
rect 8284 5866 8298 5894
rect 8138 5110 8298 5866
rect 8138 5082 8152 5110
rect 8180 5082 8204 5110
rect 8232 5082 8256 5110
rect 8284 5082 8298 5110
rect 8138 4326 8298 5082
rect 8138 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8298 4326
rect 8138 3542 8298 4298
rect 8138 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8298 3542
rect 8138 2758 8298 3514
rect 8138 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8298 2758
rect 8138 1974 8298 2730
rect 8138 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8298 1974
rect 8138 1538 8298 1946
rect 9216 7854 9376 8262
rect 9216 7826 9230 7854
rect 9258 7826 9282 7854
rect 9310 7826 9334 7854
rect 9362 7826 9376 7854
rect 9216 7070 9376 7826
rect 9216 7042 9230 7070
rect 9258 7042 9282 7070
rect 9310 7042 9334 7070
rect 9362 7042 9376 7070
rect 9216 6286 9376 7042
rect 9216 6258 9230 6286
rect 9258 6258 9282 6286
rect 9310 6258 9334 6286
rect 9362 6258 9376 6286
rect 9216 5502 9376 6258
rect 9216 5474 9230 5502
rect 9258 5474 9282 5502
rect 9310 5474 9334 5502
rect 9362 5474 9376 5502
rect 9216 4718 9376 5474
rect 9216 4690 9230 4718
rect 9258 4690 9282 4718
rect 9310 4690 9334 4718
rect 9362 4690 9376 4718
rect 9216 3934 9376 4690
rect 9216 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9376 3934
rect 9216 3150 9376 3906
rect 9216 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9376 3150
rect 9216 2366 9376 3122
rect 9216 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9376 2366
rect 9216 1582 9376 2338
rect 9216 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9376 1582
rect 9216 1538 9376 1554
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 7056
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5824 0 1 3920
box -43 -43 1051 435
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5040 0 1 7056
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5208 0 -1 3920
box -43 -43 2059 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8848 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3528 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7336 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2968 0 1 3136
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1232 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 1624 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5376 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3640 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3528 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3304 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3640 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3472 0 -1 3136
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _112_
timestamp 1698431365
transform -1 0 7056 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698431365
transform 1 0 7056 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3976 0 1 3136
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698431365
transform 1 0 7112 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 -1 3136
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _117_
timestamp 1698431365
transform -1 0 3192 0 1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698431365
transform -1 0 4704 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3864 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _120_
timestamp 1698431365
transform -1 0 2968 0 -1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3584 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2912 0 -1 4704
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698431365
transform 1 0 6720 0 1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _124_
timestamp 1698431365
transform 1 0 2968 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _125_
timestamp 1698431365
transform -1 0 6496 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _126_
timestamp 1698431365
transform 1 0 6216 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698431365
transform -1 0 6496 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1698431365
transform -1 0 4872 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3864 0 -1 5488
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698431365
transform 1 0 3920 0 -1 6272
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698431365
transform 1 0 4704 0 -1 4704
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698431365
transform 1 0 5488 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1698431365
transform -1 0 6160 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1698431365
transform -1 0 6160 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _135_
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698431365
transform 1 0 3864 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3864 0 1 6272
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4200 0 -1 6272
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1698431365
transform 1 0 6104 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698431365
transform 1 0 6160 0 -1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698431365
transform -1 0 7000 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _142_
timestamp 1698431365
transform 1 0 4816 0 1 5488
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _143_
timestamp 1698431365
transform 1 0 6048 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _144_
timestamp 1698431365
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _145_
timestamp 1698431365
transform 1 0 6384 0 -1 7056
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5488 0 1 6272
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1698431365
transform 1 0 5824 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _148_
timestamp 1698431365
transform 1 0 5040 0 -1 4704
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _149_
timestamp 1698431365
transform 1 0 4200 0 -1 7056
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5824 0 1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1698431365
transform 1 0 6888 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _152_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5768 0 -1 7056
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698431365
transform 1 0 4704 0 -1 5488
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6328 0 1 7056
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_
timestamp 1698431365
transform 1 0 5040 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _156_
timestamp 1698431365
transform -1 0 6104 0 1 6272
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698431365
transform -1 0 5824 0 1 5488
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _158_
timestamp 1698431365
transform 1 0 5880 0 1 4704
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3640 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _160_
timestamp 1698431365
transform 1 0 4816 0 -1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1698431365
transform 1 0 1344 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _162_
timestamp 1698431365
transform 1 0 1680 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _163_
timestamp 1698431365
transform 1 0 1232 0 1 3920
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698431365
transform -1 0 1792 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _165_
timestamp 1698431365
transform 1 0 1792 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _166_
timestamp 1698431365
transform 1 0 1232 0 -1 5488
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _167_
timestamp 1698431365
transform 1 0 952 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _168_
timestamp 1698431365
transform 1 0 2128 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698431365
transform -1 0 6776 0 1 1568
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698431365
transform -1 0 5376 0 -1 2352
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _171_
timestamp 1698431365
transform 1 0 6664 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _172_
timestamp 1698431365
transform -1 0 7224 0 1 2352
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _173_
timestamp 1698431365
transform 1 0 7224 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698431365
transform 1 0 7224 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698431365
transform 1 0 8904 0 -1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _176_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6664 0 1 3136
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _177_
timestamp 1698431365
transform 1 0 7224 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698431365
transform 1 0 7784 0 -1 5488
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _179_
timestamp 1698431365
transform 1 0 8008 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698431365
transform 1 0 8624 0 -1 5488
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698431365
transform -1 0 7056 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _182_
timestamp 1698431365
transform 1 0 8624 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698431365
transform 1 0 8624 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _184_
timestamp 1698431365
transform 1 0 6944 0 1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _185_
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _186_
timestamp 1698431365
transform 1 0 7000 0 1 5488
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698431365
transform 1 0 8624 0 -1 3920
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698431365
transform 1 0 8064 0 -1 5488
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _189_
timestamp 1698431365
transform 1 0 8624 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _190_
timestamp 1698431365
transform 1 0 8624 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4536 0 1 3136
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698431365
transform 1 0 2016 0 -1 2352
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698431365
transform 1 0 2744 0 1 5488
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698431365
transform 1 0 2912 0 -1 4704
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698431365
transform 1 0 2520 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698431365
transform 1 0 1848 0 -1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698431365
transform -1 0 7000 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698431365
transform 1 0 2968 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698431365
transform -1 0 7056 0 -1 3136
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698431365
transform -1 0 6496 0 1 2352
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698431365
transform 1 0 1008 0 -1 4704
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698431365
transform 1 0 1008 0 1 4704
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698431365
transform 1 0 1064 0 -1 3136
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698431365
transform 1 0 7560 0 1 3136
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698431365
transform 1 0 7560 0 1 3920
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698431365
transform 1 0 7560 0 1 5488
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698431365
transform 1 0 7560 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698431365
transform 1 0 7504 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698431365
transform 1 0 7448 0 1 4704
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8960 0 1 2352
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__A1
timestamp 1698431365
transform 1 0 2968 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__B
timestamp 1698431365
transform 1 0 9016 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__B
timestamp 1698431365
transform 1 0 9072 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698431365
transform 1 0 4424 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698431365
transform -1 0 3752 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698431365
transform 1 0 4536 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698431365
transform 1 0 4312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698431365
transform 1 0 3584 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698431365
transform -1 0 4928 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698431365
transform 1 0 2856 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698431365
transform 1 0 2520 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698431365
transform 1 0 2800 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 4816 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1232 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 1232 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 896 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 8848 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4984 0 -1 5488
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 5880 0 1 4704
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform 1 0 5712 0 -1 4704
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_28 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_32 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_52 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3584 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_55 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3752 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_63
timestamp 1698431365
transform 1 0 4200 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 4424 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_70
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_74
timestamp 1698431365
transform 1 0 4816 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_109
timestamp 1698431365
transform 1 0 6776 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138
timestamp 1698431365
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698431365
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2
timestamp 1698431365
transform 1 0 784 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_18
timestamp 1698431365
transform 1 0 1680 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_22
timestamp 1698431365
transform 1 0 1904 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_61
timestamp 1698431365
transform 1 0 4088 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 4536 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_72
timestamp 1698431365
transform 1 0 4704 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_76
timestamp 1698431365
transform 1 0 4928 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_78
timestamp 1698431365
transform 1 0 5040 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_90
timestamp 1698431365
transform 1 0 5712 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_92
timestamp 1698431365
transform 1 0 5824 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_119
timestamp 1698431365
transform 1 0 7336 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_135
timestamp 1698431365
transform 1 0 8232 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 8456 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_146
timestamp 1698431365
transform 1 0 8848 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_150
timestamp 1698431365
transform 1 0 9072 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_2
timestamp 1698431365
transform 1 0 784 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_18
timestamp 1698431365
transform 1 0 1680 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_26
timestamp 1698431365
transform 1 0 2128 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_30
timestamp 1698431365
transform 1 0 2352 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_32
timestamp 1698431365
transform 1 0 2464 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 2744 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 6496 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_107
timestamp 1698431365
transform 1 0 6664 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_148
timestamp 1698431365
transform 1 0 8960 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_2
timestamp 1698431365
transform 1 0 784 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_6
timestamp 1698431365
transform 1 0 1008 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_36
timestamp 1698431365
transform 1 0 2688 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_49
timestamp 1698431365
transform 1 0 3416 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_64
timestamp 1698431365
transform 1 0 4256 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_66
timestamp 1698431365
transform 1 0 4368 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 4536 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 4704 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_84
timestamp 1698431365
transform 1 0 5376 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 9072 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_2
timestamp 1698431365
transform 1 0 784 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_18
timestamp 1698431365
transform 1 0 1680 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_37
timestamp 1698431365
transform 1 0 2744 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_56
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_58
timestamp 1698431365
transform 1 0 3920 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_98
timestamp 1698431365
transform 1 0 6160 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 784 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_4
timestamp 1698431365
transform 1 0 896 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_17
timestamp 1698431365
transform 1 0 1624 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_34
timestamp 1698431365
transform 1 0 2576 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_38
timestamp 1698431365
transform 1 0 2800 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_40
timestamp 1698431365
transform 1 0 2912 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_61
timestamp 1698431365
transform 1 0 4088 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 4536 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_72
timestamp 1698431365
transform 1 0 4704 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_80
timestamp 1698431365
transform 1 0 5152 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_123
timestamp 1698431365
transform 1 0 7560 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 8456 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698431365
transform 1 0 1120 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 2240 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 2464 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 2744 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_41
timestamp 1698431365
transform 1 0 2968 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_49
timestamp 1698431365
transform 1 0 3416 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_51
timestamp 1698431365
transform 1 0 3528 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_60
timestamp 1698431365
transform 1 0 4032 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_68
timestamp 1698431365
transform 1 0 4480 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_71
timestamp 1698431365
transform 1 0 4648 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_73
timestamp 1698431365
transform 1 0 4760 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_96
timestamp 1698431365
transform 1 0 6048 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 6496 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_121
timestamp 1698431365
transform 1 0 7448 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_2
timestamp 1698431365
transform 1 0 784 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 4536 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_77
timestamp 1698431365
transform 1 0 4984 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_150
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698431365
transform 1 0 784 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 2744 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698431365
transform 1 0 6440 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 6664 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_120
timestamp 1698431365
transform 1 0 7392 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_150
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_2
timestamp 1698431365
transform 1 0 784 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_20
timestamp 1698431365
transform 1 0 1792 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_28
timestamp 1698431365
transform 1 0 2240 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_32
timestamp 1698431365
transform 1 0 2464 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 8344 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 8456 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_147
timestamp 1698431365
transform 1 0 8904 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_151
timestamp 1698431365
transform 1 0 9128 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_2
timestamp 1698431365
transform 1 0 784 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_10
timestamp 1698431365
transform 1 0 1232 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_20
timestamp 1698431365
transform 1 0 1792 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698431365
transform 1 0 2240 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 2464 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_72
timestamp 1698431365
transform 1 0 4704 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_84
timestamp 1698431365
transform 1 0 5376 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 6496 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 784 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_18
timestamp 1698431365
transform 1 0 1680 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_20
timestamp 1698431365
transform 1 0 1792 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_50
timestamp 1698431365
transform 1 0 3472 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_54
timestamp 1698431365
transform 1 0 3696 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 4704 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_104
timestamp 1698431365
transform 1 0 6496 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 1120 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 2240 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_37
timestamp 1698431365
transform 1 0 2744 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_53
timestamp 1698431365
transform 1 0 3640 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_75
timestamp 1698431365
transform 1 0 4872 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_103
timestamp 1698431365
transform 1 0 6440 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_107
timestamp 1698431365
transform 1 0 6664 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 784 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_18
timestamp 1698431365
transform 1 0 1680 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_26
timestamp 1698431365
transform 1 0 2128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_30
timestamp 1698431365
transform 1 0 2352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_32
timestamp 1698431365
transform 1 0 2464 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_62
timestamp 1698431365
transform 1 0 4144 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_86
timestamp 1698431365
transform 1 0 5488 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_90
timestamp 1698431365
transform 1 0 5712 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_148
timestamp 1698431365
transform 1 0 8960 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 2744 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_53
timestamp 1698431365
transform 1 0 3640 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_63
timestamp 1698431365
transform 1 0 4200 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 6664 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_111
timestamp 1698431365
transform 1 0 6888 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_151
timestamp 1698431365
transform 1 0 9128 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698431365
transform 1 0 784 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_34
timestamp 1698431365
transform 1 0 2576 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_38
timestamp 1698431365
transform 1 0 2800 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_40
timestamp 1698431365
transform 1 0 2912 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_76
timestamp 1698431365
transform 1 0 4928 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_113
timestamp 1698431365
transform 1 0 7000 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_148
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 1120 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_12
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_36
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_70
timestamp 1698431365
transform 1 0 4592 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_86
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_94
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_104
timestamp 1698431365
transform 1 0 6496 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_108
timestamp 1698431365
transform 1 0 6720 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_144
timestamp 1698431365
transform 1 0 8736 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_148
timestamp 1698431365
transform 1 0 8960 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 8736 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 784 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 784 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 784 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 9184 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2240 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698431365
transform 1 0 6832 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698431365
transform -1 0 8512 0 -1 3136
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698431365
transform -1 0 8512 0 -1 6272
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform -1 0 8512 0 -1 7056
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform -1 0 8288 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698431365
transform -1 0 8512 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform 1 0 4928 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_17 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 9296 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_18
timestamp 1698431365
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_19
timestamp 1698431365
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 9296 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_20
timestamp 1698431365
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 9296 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_21
timestamp 1698431365
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 9296 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_22
timestamp 1698431365
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 9296 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_23
timestamp 1698431365
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 9296 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_24
timestamp 1698431365
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 9296 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_25
timestamp 1698431365
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 9296 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_26
timestamp 1698431365
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 9296 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_27
timestamp 1698431365
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 9296 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_28
timestamp 1698431365
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 9296 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_29
timestamp 1698431365
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 9296 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_30
timestamp 1698431365
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 9296 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_31
timestamp 1698431365
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 9296 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_32
timestamp 1698431365
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 9296 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_33
timestamp 1698431365
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 9296 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1698431365
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_38
timestamp 1698431365
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1698431365
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_40
timestamp 1698431365
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_41
timestamp 1698431365
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_42
timestamp 1698431365
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_43
timestamp 1698431365
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_44
timestamp 1698431365
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_45
timestamp 1698431365
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_46
timestamp 1698431365
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_47
timestamp 1698431365
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_48
timestamp 1698431365
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_49
timestamp 1698431365
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_50
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_51
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_52
timestamp 1698431365
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_53
timestamp 1698431365
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_54
timestamp 1698431365
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_55
timestamp 1698431365
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_56
timestamp 1698431365
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_57
timestamp 1698431365
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_58
timestamp 1698431365
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_59
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_60
timestamp 1698431365
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_61
timestamp 1698431365
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_62
timestamp 1698431365
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_63
timestamp 1698431365
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_64
timestamp 1698431365
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_65
timestamp 1698431365
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_66
timestamp 1698431365
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_67
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_68
timestamp 1698431365
transform 1 0 2576 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_69
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_70
timestamp 1698431365
transform 1 0 6384 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_71
timestamp 1698431365
transform 1 0 8288 0 1 7840
box -43 -43 155 435
<< labels >>
flabel metal2 s 2464 9600 2520 10000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 7392 9600 7448 10000 0 FreeSans 224 90 0 0 reset
port 1 nsew signal input
flabel metal3 s 0 6160 400 6216 0 FreeSans 224 0 0 0 rle1__input_r[0]
port 2 nsew signal input
flabel metal3 s 0 8624 400 8680 0 FreeSans 224 0 0 0 rle1__input_r[1]
port 3 nsew signal input
flabel metal3 s 0 1232 400 1288 0 FreeSans 224 0 0 0 rle1__input_r_rdy
port 4 nsew signal tristate
flabel metal3 s 0 3696 400 3752 0 FreeSans 224 0 0 0 rle1__input_r_vld
port 5 nsew signal input
flabel metal3 s 9600 3024 10000 3080 0 FreeSans 224 0 0 0 rle1__output_s[0]
port 6 nsew signal tristate
flabel metal3 s 9600 4256 10000 4312 0 FreeSans 224 0 0 0 rle1__output_s[1]
port 7 nsew signal tristate
flabel metal3 s 9600 5488 10000 5544 0 FreeSans 224 0 0 0 rle1__output_s[2]
port 8 nsew signal tristate
flabel metal3 s 9600 6720 10000 6776 0 FreeSans 224 0 0 0 rle1__output_s[3]
port 9 nsew signal tristate
flabel metal3 s 9600 7952 10000 8008 0 FreeSans 224 0 0 0 rle1__output_s[4]
port 10 nsew signal tristate
flabel metal3 s 9600 9184 10000 9240 0 FreeSans 224 0 0 0 rle1__output_s[5]
port 11 nsew signal tristate
flabel metal3 s 9600 560 10000 616 0 FreeSans 224 0 0 0 rle1__output_s_rdy
port 12 nsew signal input
flabel metal3 s 9600 1792 10000 1848 0 FreeSans 224 0 0 0 rle1__output_s_vld
port 13 nsew signal tristate
flabel metal4 s 1670 1538 1830 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 3826 1538 3986 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 5982 1538 6142 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 8138 1538 8298 8262 0 FreeSans 640 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 2748 1538 2908 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 4904 1538 5064 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 7060 1538 7220 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 9216 1538 9376 8262 0 FreeSans 640 90 0 0 vss
port 15 nsew ground bidirectional
rlabel metal1 4984 8232 4984 8232 0 vdd
rlabel via1 5024 7840 5024 7840 0 vss
rlabel metal2 4228 3248 4228 3248 0 _000_
rlabel metal2 2492 2408 2492 2408 0 _001_
rlabel metal2 2884 5404 2884 5404 0 _002_
rlabel metal2 3332 4564 3332 4564 0 _003_
rlabel metal3 4116 6804 4116 6804 0 _004_
rlabel metal2 2324 5992 2324 5992 0 _005_
rlabel metal2 6216 7588 6216 7588 0 _006_
rlabel metal3 4620 7644 4620 7644 0 _007_
rlabel metal2 6580 3892 6580 3892 0 _008_
rlabel metal3 5516 2604 5516 2604 0 _009_
rlabel metal2 1484 4228 1484 4228 0 _010_
rlabel metal2 1484 5180 1484 5180 0 _011_
rlabel metal2 1540 3192 1540 3192 0 _012_
rlabel metal2 7532 3472 7532 3472 0 _013_
rlabel metal2 8148 3948 8148 3948 0 _014_
rlabel metal2 8036 5880 8036 5880 0 _015_
rlabel metal2 7420 6832 7420 6832 0 _016_
rlabel metal2 7504 5572 7504 5572 0 _017_
rlabel metal2 8764 4732 8764 4732 0 _018_
rlabel metal2 8484 2660 8484 2660 0 _019_
rlabel metal2 5600 4564 5600 4564 0 _020_
rlabel metal2 4592 6972 4592 6972 0 _021_
rlabel metal3 5908 6860 5908 6860 0 _022_
rlabel metal3 7252 6356 7252 6356 0 _023_
rlabel metal3 5096 5292 5096 5292 0 _024_
rlabel metal2 5908 6720 5908 6720 0 _025_
rlabel metal3 5180 7084 5180 7084 0 _026_
rlabel metal2 6244 5180 6244 5180 0 _027_
rlabel metal2 4032 2212 4032 2212 0 _028_
rlabel metal2 1400 4116 1400 4116 0 _029_
rlabel metal2 1596 4214 1596 4214 0 _030_
rlabel metal2 1428 5460 1428 5460 0 _031_
rlabel metal2 1596 4956 1596 4956 0 _032_
rlabel metal3 1708 3724 1708 3724 0 _033_
rlabel metal2 8876 2604 8876 2604 0 _034_
rlabel metal2 6804 2856 6804 2856 0 _035_
rlabel metal2 7364 3416 7364 3416 0 _036_
rlabel metal2 6972 2688 6972 2688 0 _037_
rlabel metal2 8652 3192 8652 3192 0 _038_
rlabel metal3 8708 3724 8708 3724 0 _039_
rlabel metal2 8708 6580 8708 6580 0 _040_
rlabel metal2 7868 5488 7868 5488 0 _041_
rlabel metal2 8008 3724 8008 3724 0 _042_
rlabel metal2 8876 5740 8876 5740 0 _043_
rlabel metal2 8652 6104 8652 6104 0 _044_
rlabel metal2 8764 7112 8764 7112 0 _045_
rlabel metal2 8820 6664 8820 6664 0 _046_
rlabel metal2 8876 4172 8876 4172 0 _047_
rlabel metal3 8540 4564 8540 4564 0 _048_
rlabel metal2 6356 2604 6356 2604 0 _049_
rlabel metal2 4284 5292 4284 5292 0 _050_
rlabel metal3 5236 4060 5236 4060 0 _051_
rlabel metal2 3948 5264 3948 5264 0 _052_
rlabel metal2 6916 3276 6916 3276 0 _053_
rlabel metal2 6692 2156 6692 2156 0 _054_
rlabel metal3 5796 2436 5796 2436 0 _055_
rlabel metal2 3948 2912 3948 2912 0 _056_
rlabel metal2 1428 3556 1428 3556 0 _057_
rlabel metal2 1596 3584 1596 3584 0 _058_
rlabel metal3 4704 3052 4704 3052 0 _059_
rlabel metal2 3332 2800 3332 2800 0 _060_
rlabel metal2 3220 3332 3220 3332 0 _061_
rlabel metal2 3808 3612 3808 3612 0 _062_
rlabel metal2 4004 3976 4004 3976 0 _063_
rlabel metal2 2828 4480 2828 4480 0 _064_
rlabel metal2 6860 5908 6860 5908 0 _065_
rlabel metal2 7308 4900 7308 4900 0 _066_
rlabel metal2 8932 3388 8932 3388 0 _067_
rlabel metal2 3136 2660 3136 2660 0 _068_
rlabel metal2 4844 4984 4844 4984 0 _069_
rlabel metal3 3304 5236 3304 5236 0 _070_
rlabel metal2 3724 4396 3724 4396 0 _071_
rlabel metal2 2660 4816 2660 4816 0 _072_
rlabel metal2 8932 5572 8932 5572 0 _073_
rlabel metal2 6328 3444 6328 3444 0 _074_
rlabel metal2 6328 5684 6328 5684 0 _075_
rlabel metal2 5180 6160 5180 6160 0 _076_
rlabel metal3 5432 6524 5432 6524 0 _077_
rlabel metal2 4452 5292 4452 5292 0 _078_
rlabel metal2 4788 4872 4788 4872 0 _079_
rlabel metal2 4788 4396 4788 4396 0 _080_
rlabel metal2 7980 5740 7980 5740 0 _081_
rlabel metal2 6076 6132 6076 6132 0 _082_
rlabel metal3 5600 5964 5600 5964 0 _083_
rlabel metal2 5292 6440 5292 6440 0 _084_
rlabel metal2 4284 6188 4284 6188 0 _085_
rlabel metal3 4732 5684 4732 5684 0 _086_
rlabel metal2 6692 7056 6692 7056 0 _087_
rlabel metal3 5740 5796 5740 5796 0 _088_
rlabel metal2 1568 4116 1568 4116 0 _089_
rlabel metal2 6356 7924 6356 7924 0 _090_
rlabel metal3 6804 7196 6804 7196 0 _091_
rlabel metal3 6356 6860 6356 6860 0 _092_
rlabel metal2 5376 6356 5376 6356 0 _093_
rlabel metal2 5936 4228 5936 4228 0 _094_
rlabel metal3 3668 6188 3668 6188 0 clk
rlabel metal2 5740 4956 5740 4956 0 clknet_0_clk
rlabel metal2 2996 7644 2996 7644 0 clknet_1_0__leaf_clk
rlabel via2 7700 2940 7700 2940 0 clknet_1_1__leaf_clk
rlabel metal2 8484 7196 8484 7196 0 net1
rlabel metal2 8904 6860 8904 6860 0 net10
rlabel metal2 8820 7896 8820 7896 0 net11
rlabel metal2 8792 3836 8792 3836 0 net12
rlabel metal3 4592 1764 4592 1764 0 net13
rlabel metal2 1428 5852 1428 5852 0 net2
rlabel metal3 1456 7924 1456 7924 0 net3
rlabel metal2 1036 3892 1036 3892 0 net4
rlabel metal2 8932 1932 8932 1932 0 net5
rlabel metal2 1260 3472 1260 3472 0 net6
rlabel metal2 7140 2576 7140 2576 0 net7
rlabel metal2 9044 3696 9044 3696 0 net8
rlabel metal2 9100 5768 9100 5768 0 net9
rlabel metal2 8596 8204 8596 8204 0 reset
rlabel metal2 868 6300 868 6300 0 rle1__input_r[0]
rlabel metal2 868 8344 868 8344 0 rle1__input_r[1]
rlabel metal3 679 1260 679 1260 0 rle1__input_r_rdy
rlabel metal3 651 3724 651 3724 0 rle1__input_r_vld
rlabel metal2 8092 2464 8092 2464 0 rle1__output_s[0]
rlabel metal2 7924 3612 7924 3612 0 rle1__output_s[1]
rlabel metal2 7924 5768 7924 5768 0 rle1__output_s[2]
rlabel metal3 8785 6748 8785 6748 0 rle1__output_s[3]
rlabel metal3 8533 7980 8533 7980 0 rle1__output_s[4]
rlabel metal2 7924 8484 7924 8484 0 rle1__output_s[5]
rlabel metal2 9100 1148 9100 1148 0 rle1__output_s_rdy
rlabel metal3 7917 1820 7917 1820 0 rle1__output_s_vld
rlabel metal2 5628 5460 5628 5460 0 rle1_enc_0.____state_0
rlabel metal2 4060 6664 4060 6664 0 rle1_enc_0.____state_1\[0\]
rlabel metal3 3668 7140 3668 7140 0 rle1_enc_0.____state_1\[1\]
rlabel metal2 5460 7784 5460 7784 0 rle1_enc_0.____state_1\[2\]
rlabel metal2 4984 7252 4984 7252 0 rle1_enc_0.____state_1\[3\]
rlabel metal2 3444 2940 3444 2940 0 rle1_enc_0.____state_2
rlabel metal2 2044 3612 2044 3612 0 rle1_enc_0.__rle1__input_r_reg\[0\]
rlabel metal3 2464 4564 2464 4564 0 rle1_enc_0.__rle1__input_r_reg\[1\]
rlabel metal2 2996 3080 2996 3080 0 rle1_enc_0.__rle1__input_r_valid_reg
rlabel metal2 6972 3416 6972 3416 0 rle1_enc_0.p0_____state_2__1
rlabel metal2 4452 4228 4452 4228 0 rle1_enc_0.p0_input_symbol
rlabel metal2 4648 5684 4648 5684 0 rle1_enc_0.p0_not_196
rlabel metal2 5236 2352 5236 2352 0 rle1_enc_0.p0_valid
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
