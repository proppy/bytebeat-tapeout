magic
tech gf180mcuD
magscale 1 10
timestamp 1702516873
<< metal1 >>
rect 48738 26798 48750 26850
rect 48802 26847 48814 26850
rect 49074 26847 49086 26850
rect 48802 26801 49086 26847
rect 48802 26798 48814 26801
rect 49074 26798 49086 26801
rect 49138 26847 49150 26850
rect 49746 26847 49758 26850
rect 49138 26801 49758 26847
rect 49138 26798 49150 26801
rect 49746 26798 49758 26801
rect 49810 26798 49822 26850
rect 1344 26682 58731 26716
rect 1344 26630 15520 26682
rect 15572 26630 15624 26682
rect 15676 26630 15728 26682
rect 15780 26630 29827 26682
rect 29879 26630 29931 26682
rect 29983 26630 30035 26682
rect 30087 26630 44134 26682
rect 44186 26630 44238 26682
rect 44290 26630 44342 26682
rect 44394 26630 58441 26682
rect 58493 26630 58545 26682
rect 58597 26630 58649 26682
rect 58701 26630 58731 26682
rect 1344 26596 58731 26630
rect 21310 26514 21362 26526
rect 12450 26462 12462 26514
rect 12514 26462 12526 26514
rect 21310 26450 21362 26462
rect 48750 26514 48802 26526
rect 48750 26450 48802 26462
rect 50318 26514 50370 26526
rect 50318 26450 50370 26462
rect 52222 26514 52274 26526
rect 52222 26450 52274 26462
rect 57710 26514 57762 26526
rect 57710 26450 57762 26462
rect 9326 26402 9378 26414
rect 20750 26402 20802 26414
rect 7970 26350 7982 26402
rect 8034 26350 8046 26402
rect 8194 26350 8206 26402
rect 8258 26350 8270 26402
rect 14018 26350 14030 26402
rect 14082 26350 14094 26402
rect 16034 26350 16046 26402
rect 16098 26350 16110 26402
rect 16370 26350 16382 26402
rect 16434 26350 16446 26402
rect 9326 26338 9378 26350
rect 20750 26338 20802 26350
rect 26686 26402 26738 26414
rect 26686 26338 26738 26350
rect 28926 26402 28978 26414
rect 49758 26402 49810 26414
rect 37426 26350 37438 26402
rect 37490 26350 37502 26402
rect 40114 26350 40126 26402
rect 40178 26350 40190 26402
rect 50642 26350 50654 26402
rect 50706 26350 50718 26402
rect 28926 26338 28978 26350
rect 49758 26338 49810 26350
rect 5518 26290 5570 26302
rect 7310 26290 7362 26302
rect 11118 26290 11170 26302
rect 22654 26290 22706 26302
rect 2146 26238 2158 26290
rect 2210 26238 2222 26290
rect 6850 26238 6862 26290
rect 6914 26238 6926 26290
rect 7186 26238 7198 26290
rect 7250 26238 7262 26290
rect 7634 26238 7646 26290
rect 7698 26238 7710 26290
rect 11330 26238 11342 26290
rect 11394 26238 11406 26290
rect 12338 26238 12350 26290
rect 12402 26238 12414 26290
rect 13234 26238 13246 26290
rect 13298 26238 13310 26290
rect 13570 26238 13582 26290
rect 13634 26238 13646 26290
rect 16258 26238 16270 26290
rect 16322 26238 16334 26290
rect 17490 26238 17502 26290
rect 17554 26238 17566 26290
rect 19170 26238 19182 26290
rect 19234 26238 19246 26290
rect 22082 26238 22094 26290
rect 22146 26238 22158 26290
rect 5518 26226 5570 26238
rect 7310 26226 7362 26238
rect 11118 26226 11170 26238
rect 22654 26226 22706 26238
rect 26910 26290 26962 26302
rect 26910 26226 26962 26238
rect 27358 26290 27410 26302
rect 29486 26290 29538 26302
rect 37998 26290 38050 26302
rect 48638 26290 48690 26302
rect 28690 26238 28702 26290
rect 28754 26238 28766 26290
rect 31266 26238 31278 26290
rect 31330 26238 31342 26290
rect 33058 26238 33070 26290
rect 33122 26238 33134 26290
rect 33730 26238 33742 26290
rect 33794 26238 33806 26290
rect 34178 26238 34190 26290
rect 34242 26238 34254 26290
rect 36194 26238 36206 26290
rect 36258 26238 36270 26290
rect 41346 26238 41358 26290
rect 41410 26238 41422 26290
rect 27358 26226 27410 26238
rect 29486 26226 29538 26238
rect 37998 26226 38050 26238
rect 48638 26226 48690 26238
rect 49534 26290 49586 26302
rect 49534 26226 49586 26238
rect 49982 26290 50034 26302
rect 49982 26226 50034 26238
rect 51326 26290 51378 26302
rect 51326 26226 51378 26238
rect 56926 26290 56978 26302
rect 56926 26226 56978 26238
rect 5070 26178 5122 26190
rect 8878 26178 8930 26190
rect 5954 26126 5966 26178
rect 6018 26126 6030 26178
rect 5070 26114 5122 26126
rect 8878 26114 8930 26126
rect 9886 26178 9938 26190
rect 20078 26178 20130 26190
rect 23102 26178 23154 26190
rect 10546 26126 10558 26178
rect 10610 26126 10622 26178
rect 19618 26126 19630 26178
rect 19682 26126 19694 26178
rect 21970 26126 21982 26178
rect 22034 26126 22046 26178
rect 9886 26114 9938 26126
rect 20078 26114 20130 26126
rect 23102 26114 23154 26126
rect 23438 26178 23490 26190
rect 23438 26114 23490 26126
rect 24670 26178 24722 26190
rect 24670 26114 24722 26126
rect 25454 26178 25506 26190
rect 25454 26114 25506 26126
rect 26014 26178 26066 26190
rect 26014 26114 26066 26126
rect 26462 26178 26514 26190
rect 26462 26114 26514 26126
rect 27134 26178 27186 26190
rect 27134 26114 27186 26126
rect 27694 26178 27746 26190
rect 32286 26178 32338 26190
rect 35422 26178 35474 26190
rect 29922 26126 29934 26178
rect 29986 26126 29998 26178
rect 33506 26126 33518 26178
rect 33570 26126 33582 26178
rect 27694 26114 27746 26126
rect 32286 26114 32338 26126
rect 35422 26114 35474 26126
rect 38558 26178 38610 26190
rect 46846 26178 46898 26190
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 38558 26114 38610 26126
rect 46846 26114 46898 26126
rect 47630 26178 47682 26190
rect 47630 26114 47682 26126
rect 48078 26178 48130 26190
rect 48078 26114 48130 26126
rect 51774 26178 51826 26190
rect 51774 26114 51826 26126
rect 53006 26178 53058 26190
rect 53006 26114 53058 26126
rect 53230 26178 53282 26190
rect 53230 26114 53282 26126
rect 56590 26178 56642 26190
rect 56590 26114 56642 26126
rect 4062 26066 4114 26078
rect 20974 26066 21026 26078
rect 15026 26014 15038 26066
rect 15090 26014 15102 26066
rect 19058 26014 19070 26066
rect 19122 26014 19134 26066
rect 4062 26002 4114 26014
rect 20974 26002 21026 26014
rect 23662 26066 23714 26078
rect 31166 26066 31218 26078
rect 42702 26066 42754 26078
rect 51214 26066 51266 26078
rect 23986 26014 23998 26066
rect 24050 26014 24062 26066
rect 29810 26014 29822 26066
rect 29874 26014 29886 26066
rect 36306 26014 36318 26066
rect 36370 26014 36382 26066
rect 49186 26014 49198 26066
rect 49250 26014 49262 26066
rect 23662 26002 23714 26014
rect 31166 26002 31218 26014
rect 42702 26002 42754 26014
rect 51214 26002 51266 26014
rect 53454 26066 53506 26078
rect 53454 26002 53506 26014
rect 53678 26066 53730 26078
rect 53678 26002 53730 26014
rect 54126 26066 54178 26078
rect 54126 26002 54178 26014
rect 1344 25898 58576 25932
rect 1344 25846 8367 25898
rect 8419 25846 8471 25898
rect 8523 25846 8575 25898
rect 8627 25846 22674 25898
rect 22726 25846 22778 25898
rect 22830 25846 22882 25898
rect 22934 25846 36981 25898
rect 37033 25846 37085 25898
rect 37137 25846 37189 25898
rect 37241 25846 51288 25898
rect 51340 25846 51392 25898
rect 51444 25846 51496 25898
rect 51548 25846 58576 25898
rect 1344 25812 58576 25846
rect 25230 25730 25282 25742
rect 37538 25678 37550 25730
rect 37602 25678 37614 25730
rect 54898 25678 54910 25730
rect 54962 25678 54974 25730
rect 25230 25666 25282 25678
rect 5854 25618 5906 25630
rect 12014 25618 12066 25630
rect 3042 25566 3054 25618
rect 3106 25566 3118 25618
rect 9762 25566 9774 25618
rect 9826 25566 9838 25618
rect 5854 25554 5906 25566
rect 12014 25554 12066 25566
rect 29374 25618 29426 25630
rect 35534 25618 35586 25630
rect 50430 25618 50482 25630
rect 30034 25566 30046 25618
rect 30098 25566 30110 25618
rect 32050 25566 32062 25618
rect 32114 25566 32126 25618
rect 42130 25566 42142 25618
rect 42194 25566 42206 25618
rect 53554 25566 53566 25618
rect 53618 25566 53630 25618
rect 29374 25554 29426 25566
rect 35534 25554 35586 25566
rect 50430 25554 50482 25566
rect 6974 25506 7026 25518
rect 1698 25454 1710 25506
rect 1762 25454 1774 25506
rect 6974 25442 7026 25454
rect 7198 25506 7250 25518
rect 11454 25506 11506 25518
rect 23102 25506 23154 25518
rect 36094 25506 36146 25518
rect 7746 25454 7758 25506
rect 7810 25454 7822 25506
rect 9426 25454 9438 25506
rect 9490 25454 9502 25506
rect 13458 25454 13470 25506
rect 13522 25454 13534 25506
rect 14354 25454 14366 25506
rect 14418 25454 14430 25506
rect 15138 25454 15150 25506
rect 15202 25454 15214 25506
rect 17154 25454 17166 25506
rect 17218 25454 17230 25506
rect 17602 25454 17614 25506
rect 17666 25454 17678 25506
rect 19730 25454 19742 25506
rect 19794 25454 19806 25506
rect 21522 25454 21534 25506
rect 21586 25454 21598 25506
rect 24658 25454 24670 25506
rect 24722 25454 24734 25506
rect 26114 25454 26126 25506
rect 26178 25454 26190 25506
rect 27682 25454 27694 25506
rect 27746 25454 27758 25506
rect 30146 25454 30158 25506
rect 30210 25454 30222 25506
rect 32386 25454 32398 25506
rect 32450 25454 32462 25506
rect 32834 25454 32846 25506
rect 32898 25454 32910 25506
rect 34514 25454 34526 25506
rect 34578 25454 34590 25506
rect 7198 25442 7250 25454
rect 11454 25442 11506 25454
rect 23102 25442 23154 25454
rect 36094 25442 36146 25454
rect 36430 25506 36482 25518
rect 36430 25442 36482 25454
rect 36990 25506 37042 25518
rect 51886 25506 51938 25518
rect 37202 25454 37214 25506
rect 37266 25454 37278 25506
rect 38770 25454 38782 25506
rect 38834 25454 38846 25506
rect 38994 25454 39006 25506
rect 39058 25454 39070 25506
rect 41794 25454 41806 25506
rect 41858 25454 41870 25506
rect 45378 25454 45390 25506
rect 45442 25454 45454 25506
rect 46498 25454 46510 25506
rect 46562 25454 46574 25506
rect 48626 25454 48638 25506
rect 48690 25454 48702 25506
rect 36990 25442 37042 25454
rect 51886 25442 51938 25454
rect 52110 25506 52162 25518
rect 53442 25454 53454 25506
rect 53506 25454 53518 25506
rect 55458 25454 55470 25506
rect 55522 25454 55534 25506
rect 52110 25442 52162 25454
rect 9102 25394 9154 25406
rect 8082 25342 8094 25394
rect 8146 25342 8158 25394
rect 9102 25330 9154 25342
rect 12910 25394 12962 25406
rect 12910 25330 12962 25342
rect 16718 25394 16770 25406
rect 23886 25394 23938 25406
rect 25566 25394 25618 25406
rect 35870 25394 35922 25406
rect 20178 25342 20190 25394
rect 20242 25342 20254 25394
rect 21298 25342 21310 25394
rect 21362 25342 21374 25394
rect 24434 25342 24446 25394
rect 24498 25342 24510 25394
rect 26674 25342 26686 25394
rect 26738 25342 26750 25394
rect 28466 25342 28478 25394
rect 28530 25342 28542 25394
rect 32722 25342 32734 25394
rect 32786 25342 32798 25394
rect 16718 25330 16770 25342
rect 23886 25330 23938 25342
rect 25566 25330 25618 25342
rect 35870 25330 35922 25342
rect 42702 25394 42754 25406
rect 49198 25394 49250 25406
rect 45154 25342 45166 25394
rect 45218 25342 45230 25394
rect 42702 25330 42754 25342
rect 49198 25330 49250 25342
rect 5182 25282 5234 25294
rect 5182 25218 5234 25230
rect 6302 25282 6354 25294
rect 12350 25282 12402 25294
rect 6626 25230 6638 25282
rect 6690 25230 6702 25282
rect 6302 25218 6354 25230
rect 12350 25218 12402 25230
rect 13582 25282 13634 25294
rect 13582 25218 13634 25230
rect 16494 25282 16546 25294
rect 16494 25218 16546 25230
rect 16606 25282 16658 25294
rect 16606 25218 16658 25230
rect 20638 25282 20690 25294
rect 20638 25218 20690 25230
rect 23326 25282 23378 25294
rect 23326 25218 23378 25230
rect 34974 25282 35026 25294
rect 34974 25218 35026 25230
rect 36318 25282 36370 25294
rect 36318 25218 36370 25230
rect 43262 25282 43314 25294
rect 43262 25218 43314 25230
rect 48190 25282 48242 25294
rect 48190 25218 48242 25230
rect 50206 25282 50258 25294
rect 52894 25282 52946 25294
rect 51538 25230 51550 25282
rect 51602 25230 51614 25282
rect 50206 25218 50258 25230
rect 52894 25218 52946 25230
rect 1344 25114 58731 25148
rect 1344 25062 15520 25114
rect 15572 25062 15624 25114
rect 15676 25062 15728 25114
rect 15780 25062 29827 25114
rect 29879 25062 29931 25114
rect 29983 25062 30035 25114
rect 30087 25062 44134 25114
rect 44186 25062 44238 25114
rect 44290 25062 44342 25114
rect 44394 25062 58441 25114
rect 58493 25062 58545 25114
rect 58597 25062 58649 25114
rect 58701 25062 58731 25114
rect 1344 25028 58731 25062
rect 9774 24946 9826 24958
rect 9774 24882 9826 24894
rect 25566 24946 25618 24958
rect 25566 24882 25618 24894
rect 31390 24946 31442 24958
rect 34078 24946 34130 24958
rect 39678 24946 39730 24958
rect 31714 24894 31726 24946
rect 31778 24894 31790 24946
rect 35858 24894 35870 24946
rect 35922 24894 35934 24946
rect 31390 24882 31442 24894
rect 34078 24882 34130 24894
rect 39678 24882 39730 24894
rect 47854 24946 47906 24958
rect 47854 24882 47906 24894
rect 49198 24946 49250 24958
rect 49198 24882 49250 24894
rect 5630 24834 5682 24846
rect 27246 24834 27298 24846
rect 8754 24782 8766 24834
rect 8818 24782 8830 24834
rect 11890 24782 11902 24834
rect 11954 24782 11966 24834
rect 12898 24782 12910 24834
rect 12962 24782 12974 24834
rect 21410 24782 21422 24834
rect 21474 24782 21486 24834
rect 22642 24782 22654 24834
rect 22706 24782 22718 24834
rect 24658 24782 24670 24834
rect 24722 24782 24734 24834
rect 5630 24770 5682 24782
rect 27246 24770 27298 24782
rect 29150 24834 29202 24846
rect 29150 24770 29202 24782
rect 32174 24834 32226 24846
rect 32174 24770 32226 24782
rect 33182 24834 33234 24846
rect 33182 24770 33234 24782
rect 33406 24834 33458 24846
rect 33406 24770 33458 24782
rect 33742 24834 33794 24846
rect 33742 24770 33794 24782
rect 33854 24834 33906 24846
rect 37438 24834 37490 24846
rect 49646 24834 49698 24846
rect 34962 24782 34974 24834
rect 35026 24782 35038 24834
rect 44706 24782 44718 24834
rect 44770 24782 44782 24834
rect 33854 24770 33906 24782
rect 37438 24770 37490 24782
rect 49646 24770 49698 24782
rect 53006 24834 53058 24846
rect 54898 24782 54910 24834
rect 54962 24782 54974 24834
rect 53006 24770 53058 24782
rect 2494 24722 2546 24734
rect 2494 24658 2546 24670
rect 3166 24722 3218 24734
rect 4958 24722 5010 24734
rect 14926 24722 14978 24734
rect 26686 24722 26738 24734
rect 3714 24670 3726 24722
rect 3778 24670 3790 24722
rect 5394 24670 5406 24722
rect 5458 24670 5470 24722
rect 6402 24670 6414 24722
rect 6466 24670 6478 24722
rect 7634 24670 7646 24722
rect 7698 24670 7710 24722
rect 10210 24670 10222 24722
rect 10274 24670 10286 24722
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 15138 24670 15150 24722
rect 15202 24670 15214 24722
rect 17490 24670 17502 24722
rect 17554 24670 17566 24722
rect 18386 24670 18398 24722
rect 18450 24670 18462 24722
rect 19058 24670 19070 24722
rect 19122 24670 19134 24722
rect 20402 24670 20414 24722
rect 20466 24670 20478 24722
rect 22530 24670 22542 24722
rect 22594 24670 22606 24722
rect 25666 24670 25678 24722
rect 25730 24670 25742 24722
rect 3166 24658 3218 24670
rect 4958 24658 5010 24670
rect 14926 24658 14978 24670
rect 26686 24658 26738 24670
rect 28366 24722 28418 24734
rect 30494 24722 30546 24734
rect 30146 24670 30158 24722
rect 30210 24670 30222 24722
rect 28366 24658 28418 24670
rect 30494 24658 30546 24670
rect 32062 24722 32114 24734
rect 38558 24722 38610 24734
rect 42366 24722 42418 24734
rect 36418 24670 36430 24722
rect 36482 24670 36494 24722
rect 39554 24670 39566 24722
rect 39618 24670 39630 24722
rect 42018 24670 42030 24722
rect 42082 24670 42094 24722
rect 32062 24658 32114 24670
rect 38558 24658 38610 24670
rect 42366 24658 42418 24670
rect 42702 24722 42754 24734
rect 43262 24722 43314 24734
rect 50878 24722 50930 24734
rect 43026 24670 43038 24722
rect 43090 24670 43102 24722
rect 45938 24670 45950 24722
rect 46002 24670 46014 24722
rect 49074 24670 49086 24722
rect 49138 24670 49150 24722
rect 52434 24670 52446 24722
rect 52498 24670 52510 24722
rect 54562 24670 54574 24722
rect 54626 24670 54638 24722
rect 42702 24658 42754 24670
rect 43262 24658 43314 24670
rect 50878 24658 50930 24670
rect 7198 24610 7250 24622
rect 9886 24610 9938 24622
rect 14590 24610 14642 24622
rect 27806 24610 27858 24622
rect 42926 24610 42978 24622
rect 48190 24610 48242 24622
rect 53454 24610 53506 24622
rect 56590 24610 56642 24622
rect 8978 24558 8990 24610
rect 9042 24558 9054 24610
rect 10434 24558 10446 24610
rect 10498 24558 10510 24610
rect 13906 24558 13918 24610
rect 13970 24558 13982 24610
rect 16146 24558 16158 24610
rect 16210 24558 16222 24610
rect 18274 24558 18286 24610
rect 18338 24558 18350 24610
rect 21186 24558 21198 24610
rect 21250 24558 21262 24610
rect 22306 24558 22318 24610
rect 22370 24558 22382 24610
rect 25778 24558 25790 24610
rect 25842 24558 25854 24610
rect 30930 24558 30942 24610
rect 30994 24558 31006 24610
rect 33058 24558 33070 24610
rect 33122 24558 33134 24610
rect 39330 24558 39342 24610
rect 39394 24558 39406 24610
rect 42242 24558 42254 24610
rect 42306 24558 42318 24610
rect 44482 24558 44494 24610
rect 44546 24558 44558 24610
rect 52098 24558 52110 24610
rect 52162 24558 52174 24610
rect 55234 24558 55246 24610
rect 55298 24558 55310 24610
rect 7198 24546 7250 24558
rect 9886 24546 9938 24558
rect 14590 24546 14642 24558
rect 27806 24546 27858 24558
rect 42926 24546 42978 24558
rect 48190 24546 48242 24558
rect 53454 24546 53506 24558
rect 56590 24546 56642 24558
rect 1710 24498 1762 24510
rect 1710 24434 1762 24446
rect 6638 24498 6690 24510
rect 6638 24434 6690 24446
rect 17502 24498 17554 24510
rect 32174 24498 32226 24510
rect 22194 24446 22206 24498
rect 22258 24446 22270 24498
rect 17502 24434 17554 24446
rect 32174 24434 32226 24446
rect 47294 24498 47346 24510
rect 56814 24498 56866 24510
rect 47506 24446 47518 24498
rect 47570 24495 47582 24498
rect 48066 24495 48078 24498
rect 47570 24449 48078 24495
rect 47570 24446 47582 24449
rect 48066 24446 48078 24449
rect 48130 24446 48142 24498
rect 57138 24446 57150 24498
rect 57202 24446 57214 24498
rect 47294 24434 47346 24446
rect 56814 24434 56866 24446
rect 1344 24330 58576 24364
rect 1344 24278 8367 24330
rect 8419 24278 8471 24330
rect 8523 24278 8575 24330
rect 8627 24278 22674 24330
rect 22726 24278 22778 24330
rect 22830 24278 22882 24330
rect 22934 24278 36981 24330
rect 37033 24278 37085 24330
rect 37137 24278 37189 24330
rect 37241 24278 51288 24330
rect 51340 24278 51392 24330
rect 51444 24278 51496 24330
rect 51548 24278 58576 24330
rect 1344 24244 58576 24278
rect 21646 24162 21698 24174
rect 21646 24098 21698 24110
rect 36094 24162 36146 24174
rect 36094 24098 36146 24110
rect 30606 24050 30658 24062
rect 3266 23998 3278 24050
rect 3330 23998 3342 24050
rect 8866 23998 8878 24050
rect 8930 23998 8942 24050
rect 12898 23998 12910 24050
rect 12962 23998 12974 24050
rect 15250 23998 15262 24050
rect 15314 23998 15326 24050
rect 20066 23998 20078 24050
rect 20130 23998 20142 24050
rect 22082 23998 22094 24050
rect 22146 23998 22158 24050
rect 30606 23986 30658 23998
rect 33630 24050 33682 24062
rect 33630 23986 33682 23998
rect 34750 24050 34802 24062
rect 35982 24050 36034 24062
rect 35298 23998 35310 24050
rect 35362 23998 35374 24050
rect 42914 23998 42926 24050
rect 42978 23998 42990 24050
rect 51090 23998 51102 24050
rect 51154 23998 51166 24050
rect 34750 23986 34802 23998
rect 35982 23986 36034 23998
rect 15710 23938 15762 23950
rect 18510 23938 18562 23950
rect 21870 23938 21922 23950
rect 46846 23938 46898 23950
rect 3042 23886 3054 23938
rect 3106 23886 3118 23938
rect 7746 23886 7758 23938
rect 7810 23886 7822 23938
rect 10322 23886 10334 23938
rect 10386 23886 10398 23938
rect 10770 23886 10782 23938
rect 10834 23886 10846 23938
rect 10994 23886 11006 23938
rect 11058 23886 11070 23938
rect 11330 23886 11342 23938
rect 11394 23886 11406 23938
rect 12226 23886 12238 23938
rect 12290 23886 12302 23938
rect 14914 23886 14926 23938
rect 14978 23886 14990 23938
rect 16146 23886 16158 23938
rect 16210 23886 16222 23938
rect 16706 23886 16718 23938
rect 16770 23886 16782 23938
rect 19954 23886 19966 23938
rect 20018 23886 20030 23938
rect 24322 23886 24334 23938
rect 24386 23886 24398 23938
rect 24770 23886 24782 23938
rect 24834 23886 24846 23938
rect 27346 23886 27358 23938
rect 27410 23886 27422 23938
rect 27794 23886 27806 23938
rect 27858 23886 27870 23938
rect 28466 23886 28478 23938
rect 28530 23886 28542 23938
rect 29138 23886 29150 23938
rect 29202 23886 29214 23938
rect 31042 23886 31054 23938
rect 31106 23886 31118 23938
rect 32834 23886 32846 23938
rect 32898 23886 32910 23938
rect 35746 23886 35758 23938
rect 35810 23886 35822 23938
rect 37874 23886 37886 23938
rect 37938 23886 37950 23938
rect 39218 23886 39230 23938
rect 39282 23886 39294 23938
rect 41010 23886 41022 23938
rect 41074 23886 41086 23938
rect 42802 23886 42814 23938
rect 42866 23886 42878 23938
rect 47170 23886 47182 23938
rect 47234 23886 47246 23938
rect 49522 23886 49534 23938
rect 49586 23886 49598 23938
rect 51538 23886 51550 23938
rect 51602 23886 51614 23938
rect 53106 23886 53118 23938
rect 53170 23886 53182 23938
rect 53554 23886 53566 23938
rect 53618 23886 53630 23938
rect 55570 23886 55582 23938
rect 55634 23886 55646 23938
rect 56578 23886 56590 23938
rect 56642 23886 56654 23938
rect 57922 23886 57934 23938
rect 57986 23886 57998 23938
rect 15710 23874 15762 23886
rect 18510 23874 18562 23886
rect 21870 23874 21922 23886
rect 46846 23874 46898 23886
rect 20526 23826 20578 23838
rect 4610 23774 4622 23826
rect 4674 23774 4686 23826
rect 5730 23774 5742 23826
rect 5794 23774 5806 23826
rect 8082 23774 8094 23826
rect 8146 23774 8158 23826
rect 9090 23774 9102 23826
rect 9154 23774 9166 23826
rect 12338 23774 12350 23826
rect 12402 23774 12414 23826
rect 18162 23774 18174 23826
rect 18226 23774 18238 23826
rect 20526 23762 20578 23774
rect 20638 23826 20690 23838
rect 20638 23762 20690 23774
rect 22206 23826 22258 23838
rect 22206 23762 22258 23774
rect 22430 23826 22482 23838
rect 25342 23826 25394 23838
rect 35086 23826 35138 23838
rect 44270 23826 44322 23838
rect 22754 23774 22766 23826
rect 22818 23774 22830 23826
rect 27906 23774 27918 23826
rect 27970 23774 27982 23826
rect 29250 23774 29262 23826
rect 29314 23774 29326 23826
rect 31714 23774 31726 23826
rect 31778 23774 31790 23826
rect 32722 23774 32734 23826
rect 32786 23774 32798 23826
rect 37538 23774 37550 23826
rect 37602 23774 37614 23826
rect 41682 23774 41694 23826
rect 41746 23774 41758 23826
rect 22430 23762 22482 23774
rect 25342 23762 25394 23774
rect 35086 23762 35138 23774
rect 44270 23762 44322 23774
rect 47070 23826 47122 23838
rect 48626 23774 48638 23826
rect 48690 23774 48702 23826
rect 49634 23774 49646 23826
rect 49698 23774 49710 23826
rect 51314 23774 51326 23826
rect 51378 23774 51390 23826
rect 54226 23774 54238 23826
rect 54290 23774 54302 23826
rect 55794 23774 55806 23826
rect 55858 23774 55870 23826
rect 47070 23762 47122 23774
rect 2270 23714 2322 23726
rect 2270 23650 2322 23662
rect 5070 23714 5122 23726
rect 12014 23714 12066 23726
rect 6626 23662 6638 23714
rect 6690 23662 6702 23714
rect 8306 23662 8318 23714
rect 8370 23662 8382 23714
rect 5070 23650 5122 23662
rect 12014 23650 12066 23662
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 20862 23714 20914 23726
rect 35310 23714 35362 23726
rect 46286 23714 46338 23726
rect 26450 23662 26462 23714
rect 26514 23662 26526 23714
rect 29698 23662 29710 23714
rect 29762 23662 29774 23714
rect 38546 23662 38558 23714
rect 38610 23662 38622 23714
rect 20862 23650 20914 23662
rect 35310 23650 35362 23662
rect 46286 23650 46338 23662
rect 52110 23714 52162 23726
rect 52110 23650 52162 23662
rect 54798 23714 54850 23726
rect 57598 23714 57650 23726
rect 56466 23662 56478 23714
rect 56530 23662 56542 23714
rect 54798 23650 54850 23662
rect 57598 23650 57650 23662
rect 1344 23546 58731 23580
rect 1344 23494 15520 23546
rect 15572 23494 15624 23546
rect 15676 23494 15728 23546
rect 15780 23494 29827 23546
rect 29879 23494 29931 23546
rect 29983 23494 30035 23546
rect 30087 23494 44134 23546
rect 44186 23494 44238 23546
rect 44290 23494 44342 23546
rect 44394 23494 58441 23546
rect 58493 23494 58545 23546
rect 58597 23494 58649 23546
rect 58701 23494 58731 23546
rect 1344 23460 58731 23494
rect 16942 23378 16994 23390
rect 16942 23314 16994 23326
rect 22318 23378 22370 23390
rect 22318 23314 22370 23326
rect 22542 23378 22594 23390
rect 22542 23314 22594 23326
rect 24558 23378 24610 23390
rect 24558 23314 24610 23326
rect 52670 23378 52722 23390
rect 52670 23314 52722 23326
rect 1710 23266 1762 23278
rect 1710 23202 1762 23214
rect 2942 23266 2994 23278
rect 24446 23266 24498 23278
rect 52110 23266 52162 23278
rect 10658 23214 10670 23266
rect 10722 23214 10734 23266
rect 13458 23214 13470 23266
rect 13522 23214 13534 23266
rect 16146 23214 16158 23266
rect 16210 23214 16222 23266
rect 28018 23214 28030 23266
rect 28082 23214 28094 23266
rect 28690 23214 28702 23266
rect 28754 23214 28766 23266
rect 35298 23214 35310 23266
rect 35362 23214 35374 23266
rect 38210 23214 38222 23266
rect 38274 23214 38286 23266
rect 47282 23214 47294 23266
rect 47346 23214 47358 23266
rect 49522 23214 49534 23266
rect 49586 23214 49598 23266
rect 50530 23214 50542 23266
rect 50594 23214 50606 23266
rect 2942 23202 2994 23214
rect 24446 23202 24498 23214
rect 52110 23202 52162 23214
rect 52446 23266 52498 23278
rect 52446 23202 52498 23214
rect 55470 23266 55522 23278
rect 55470 23202 55522 23214
rect 22654 23154 22706 23166
rect 23886 23154 23938 23166
rect 2482 23102 2494 23154
rect 2546 23102 2558 23154
rect 3714 23102 3726 23154
rect 3778 23102 3790 23154
rect 5954 23102 5966 23154
rect 6018 23102 6030 23154
rect 6738 23102 6750 23154
rect 6802 23102 6814 23154
rect 8754 23102 8766 23154
rect 8818 23102 8830 23154
rect 9762 23102 9774 23154
rect 9826 23102 9838 23154
rect 11442 23102 11454 23154
rect 11506 23102 11518 23154
rect 12674 23102 12686 23154
rect 12738 23102 12750 23154
rect 14466 23102 14478 23154
rect 14530 23102 14542 23154
rect 16482 23102 16494 23154
rect 16546 23102 16558 23154
rect 18274 23102 18286 23154
rect 18338 23102 18350 23154
rect 19954 23102 19966 23154
rect 20018 23102 20030 23154
rect 21970 23102 21982 23154
rect 22034 23102 22046 23154
rect 23314 23102 23326 23154
rect 23378 23102 23390 23154
rect 22654 23090 22706 23102
rect 23886 23090 23938 23102
rect 24782 23154 24834 23166
rect 24782 23090 24834 23102
rect 25230 23154 25282 23166
rect 37102 23154 37154 23166
rect 27122 23102 27134 23154
rect 27186 23102 27198 23154
rect 30370 23102 30382 23154
rect 30434 23102 30446 23154
rect 30818 23102 30830 23154
rect 30882 23102 30894 23154
rect 31042 23102 31054 23154
rect 31106 23102 31118 23154
rect 32050 23102 32062 23154
rect 32114 23102 32126 23154
rect 33730 23102 33742 23154
rect 33794 23102 33806 23154
rect 35410 23102 35422 23154
rect 35474 23102 35486 23154
rect 36866 23102 36878 23154
rect 36930 23102 36942 23154
rect 25230 23090 25282 23102
rect 37102 23090 37154 23102
rect 40350 23154 40402 23166
rect 42254 23154 42306 23166
rect 51886 23154 51938 23166
rect 41234 23102 41246 23154
rect 41298 23102 41310 23154
rect 41570 23102 41582 23154
rect 41634 23102 41646 23154
rect 42914 23102 42926 23154
rect 42978 23102 42990 23154
rect 46498 23102 46510 23154
rect 46562 23102 46574 23154
rect 47058 23102 47070 23154
rect 47122 23102 47134 23154
rect 48738 23102 48750 23154
rect 48802 23102 48814 23154
rect 40350 23090 40402 23102
rect 42254 23090 42306 23102
rect 51886 23090 51938 23102
rect 52334 23154 52386 23166
rect 52334 23090 52386 23102
rect 53454 23154 53506 23166
rect 53454 23090 53506 23102
rect 53678 23154 53730 23166
rect 53678 23090 53730 23102
rect 54126 23154 54178 23166
rect 54786 23102 54798 23154
rect 54850 23102 54862 23154
rect 56914 23102 56926 23154
rect 56978 23102 56990 23154
rect 54126 23090 54178 23102
rect 2718 23042 2770 23054
rect 17614 23042 17666 23054
rect 21086 23042 21138 23054
rect 26462 23042 26514 23054
rect 36318 23042 36370 23054
rect 53006 23042 53058 23054
rect 3602 22990 3614 23042
rect 3666 22990 3678 23042
rect 6290 22990 6302 23042
rect 6354 22990 6366 23042
rect 8082 22990 8094 23042
rect 8146 22990 8158 23042
rect 11666 22990 11678 23042
rect 11730 22990 11742 23042
rect 17826 22990 17838 23042
rect 17890 22990 17902 23042
rect 19730 22990 19742 23042
rect 19794 22990 19806 23042
rect 23426 22990 23438 23042
rect 23490 22990 23502 23042
rect 25666 22990 25678 23042
rect 25730 22990 25742 23042
rect 26786 22990 26798 23042
rect 26850 22990 26862 23042
rect 30482 22990 30494 23042
rect 30546 22990 30558 23042
rect 33618 22990 33630 23042
rect 33682 22990 33694 23042
rect 34738 22990 34750 23042
rect 34802 22990 34814 23042
rect 37650 22990 37662 23042
rect 37714 22990 37726 23042
rect 39890 22990 39902 23042
rect 39954 22990 39966 23042
rect 41346 22990 41358 23042
rect 41410 22990 41422 23042
rect 43026 22990 43038 23042
rect 43090 22990 43102 23042
rect 44594 22990 44606 23042
rect 44658 22990 44670 23042
rect 46946 22990 46958 23042
rect 47010 22990 47022 23042
rect 2718 22978 2770 22990
rect 17614 22978 17666 22990
rect 21086 22978 21138 22990
rect 26462 22978 26514 22990
rect 36318 22978 36370 22990
rect 53006 22978 53058 22990
rect 53566 23042 53618 23054
rect 55918 23042 55970 23054
rect 54674 22990 54686 23042
rect 54738 22990 54750 23042
rect 57026 22990 57038 23042
rect 57090 22990 57102 23042
rect 53566 22978 53618 22990
rect 55918 22978 55970 22990
rect 1822 22930 1874 22942
rect 35982 22930 36034 22942
rect 4834 22878 4846 22930
rect 4898 22878 4910 22930
rect 31266 22878 31278 22930
rect 31330 22878 31342 22930
rect 1822 22866 1874 22878
rect 35982 22866 36034 22878
rect 37214 22930 37266 22942
rect 37214 22866 37266 22878
rect 39006 22930 39058 22942
rect 57250 22878 57262 22930
rect 57314 22878 57326 22930
rect 39006 22866 39058 22878
rect 1344 22762 58576 22796
rect 1344 22710 8367 22762
rect 8419 22710 8471 22762
rect 8523 22710 8575 22762
rect 8627 22710 22674 22762
rect 22726 22710 22778 22762
rect 22830 22710 22882 22762
rect 22934 22710 36981 22762
rect 37033 22710 37085 22762
rect 37137 22710 37189 22762
rect 37241 22710 51288 22762
rect 51340 22710 51392 22762
rect 51444 22710 51496 22762
rect 51548 22710 58576 22762
rect 1344 22676 58576 22710
rect 24670 22594 24722 22606
rect 35198 22594 35250 22606
rect 51662 22594 51714 22606
rect 11890 22542 11902 22594
rect 11954 22542 11966 22594
rect 27122 22542 27134 22594
rect 27186 22542 27198 22594
rect 49410 22542 49422 22594
rect 49474 22542 49486 22594
rect 24670 22530 24722 22542
rect 35198 22530 35250 22542
rect 51662 22530 51714 22542
rect 10770 22430 10782 22482
rect 10834 22430 10846 22482
rect 20178 22430 20190 22482
rect 20242 22430 20254 22482
rect 22194 22430 22206 22482
rect 22258 22430 22270 22482
rect 38098 22430 38110 22482
rect 38162 22430 38174 22482
rect 40338 22430 40350 22482
rect 40402 22430 40414 22482
rect 41458 22430 41470 22482
rect 41522 22430 41534 22482
rect 44258 22430 44270 22482
rect 44322 22430 44334 22482
rect 8542 22370 8594 22382
rect 2370 22318 2382 22370
rect 2434 22318 2446 22370
rect 4386 22318 4398 22370
rect 4450 22318 4462 22370
rect 7186 22318 7198 22370
rect 7250 22318 7262 22370
rect 7746 22318 7758 22370
rect 7810 22318 7822 22370
rect 8542 22306 8594 22318
rect 8878 22370 8930 22382
rect 13582 22370 13634 22382
rect 17838 22370 17890 22382
rect 20414 22370 20466 22382
rect 24334 22370 24386 22382
rect 9090 22318 9102 22370
rect 9154 22318 9166 22370
rect 10882 22318 10894 22370
rect 10946 22318 10958 22370
rect 15250 22318 15262 22370
rect 15314 22318 15326 22370
rect 17266 22318 17278 22370
rect 17330 22318 17342 22370
rect 18610 22318 18622 22370
rect 18674 22318 18686 22370
rect 21522 22318 21534 22370
rect 21586 22318 21598 22370
rect 22978 22318 22990 22370
rect 23042 22318 23054 22370
rect 8878 22306 8930 22318
rect 13582 22306 13634 22318
rect 17838 22306 17890 22318
rect 20414 22306 20466 22318
rect 24334 22306 24386 22318
rect 26574 22370 26626 22382
rect 51438 22370 51490 22382
rect 27122 22318 27134 22370
rect 27186 22318 27198 22370
rect 29586 22318 29598 22370
rect 29650 22318 29662 22370
rect 30146 22318 30158 22370
rect 30210 22318 30222 22370
rect 32050 22318 32062 22370
rect 32114 22318 32126 22370
rect 32722 22318 32734 22370
rect 32786 22318 32798 22370
rect 33506 22318 33518 22370
rect 33570 22318 33582 22370
rect 38210 22318 38222 22370
rect 38274 22318 38286 22370
rect 40002 22318 40014 22370
rect 40066 22318 40078 22370
rect 41010 22318 41022 22370
rect 41074 22318 41086 22370
rect 43586 22318 43598 22370
rect 43650 22318 43662 22370
rect 45938 22318 45950 22370
rect 46002 22318 46014 22370
rect 47058 22318 47070 22370
rect 47122 22318 47134 22370
rect 48402 22318 48414 22370
rect 48466 22318 48478 22370
rect 49522 22318 49534 22370
rect 49586 22318 49598 22370
rect 50642 22318 50654 22370
rect 50706 22318 50718 22370
rect 26574 22306 26626 22318
rect 51438 22306 51490 22318
rect 52782 22370 52834 22382
rect 52782 22306 52834 22318
rect 53006 22370 53058 22382
rect 54338 22318 54350 22370
rect 54402 22318 54414 22370
rect 56354 22318 56366 22370
rect 56418 22318 56430 22370
rect 53006 22306 53058 22318
rect 8206 22258 8258 22270
rect 20750 22258 20802 22270
rect 2706 22206 2718 22258
rect 2770 22206 2782 22258
rect 4610 22206 4622 22258
rect 4674 22206 4686 22258
rect 6178 22206 6190 22258
rect 6242 22206 6254 22258
rect 13682 22206 13694 22258
rect 13746 22206 13758 22258
rect 14242 22206 14254 22258
rect 14306 22206 14318 22258
rect 15922 22206 15934 22258
rect 15986 22206 15998 22258
rect 8206 22194 8258 22206
rect 20750 22194 20802 22206
rect 22430 22258 22482 22270
rect 26798 22258 26850 22270
rect 53230 22258 53282 22270
rect 23538 22206 23550 22258
rect 23602 22206 23614 22258
rect 23986 22206 23998 22258
rect 24050 22206 24062 22258
rect 25666 22206 25678 22258
rect 25730 22206 25742 22258
rect 26226 22206 26238 22258
rect 26290 22206 26302 22258
rect 28242 22206 28254 22258
rect 28306 22206 28318 22258
rect 30818 22206 30830 22258
rect 30882 22206 30894 22258
rect 33394 22206 33406 22258
rect 33458 22206 33470 22258
rect 34402 22206 34414 22258
rect 34466 22206 34478 22258
rect 34850 22206 34862 22258
rect 34914 22206 34926 22258
rect 44034 22206 44046 22258
rect 44098 22206 44110 22258
rect 46050 22206 46062 22258
rect 46114 22206 46126 22258
rect 47954 22206 47966 22258
rect 48018 22206 48030 22258
rect 22430 22194 22482 22206
rect 26798 22194 26850 22206
rect 53230 22194 53282 22206
rect 53678 22258 53730 22270
rect 53678 22194 53730 22206
rect 53790 22258 53842 22270
rect 53790 22194 53842 22206
rect 55470 22258 55522 22270
rect 55470 22194 55522 22206
rect 57486 22258 57538 22270
rect 57486 22194 57538 22206
rect 8318 22146 8370 22158
rect 3378 22094 3390 22146
rect 3442 22094 3454 22146
rect 8318 22082 8370 22094
rect 13022 22146 13074 22158
rect 15038 22146 15090 22158
rect 13794 22094 13806 22146
rect 13858 22094 13870 22146
rect 13022 22082 13074 22094
rect 15038 22082 15090 22094
rect 22766 22146 22818 22158
rect 22766 22082 22818 22094
rect 25342 22146 25394 22158
rect 25342 22082 25394 22094
rect 35534 22146 35586 22158
rect 52894 22146 52946 22158
rect 46946 22094 46958 22146
rect 47010 22094 47022 22146
rect 51986 22094 51998 22146
rect 52050 22094 52062 22146
rect 35534 22082 35586 22094
rect 52894 22082 52946 22094
rect 54014 22146 54066 22158
rect 56466 22094 56478 22146
rect 56530 22094 56542 22146
rect 54014 22082 54066 22094
rect 1344 21978 58731 22012
rect 1344 21926 15520 21978
rect 15572 21926 15624 21978
rect 15676 21926 15728 21978
rect 15780 21926 29827 21978
rect 29879 21926 29931 21978
rect 29983 21926 30035 21978
rect 30087 21926 44134 21978
rect 44186 21926 44238 21978
rect 44290 21926 44342 21978
rect 44394 21926 58441 21978
rect 58493 21926 58545 21978
rect 58597 21926 58649 21978
rect 58701 21926 58731 21978
rect 1344 21892 58731 21926
rect 3390 21810 3442 21822
rect 17726 21810 17778 21822
rect 8866 21758 8878 21810
rect 8930 21758 8942 21810
rect 12786 21758 12798 21810
rect 12850 21758 12862 21810
rect 3390 21746 3442 21758
rect 17726 21746 17778 21758
rect 22766 21810 22818 21822
rect 52334 21810 52386 21822
rect 26562 21758 26574 21810
rect 26626 21758 26638 21810
rect 54226 21758 54238 21810
rect 54290 21758 54302 21810
rect 22766 21746 22818 21758
rect 52334 21746 52386 21758
rect 14366 21698 14418 21710
rect 24558 21698 24610 21710
rect 42142 21698 42194 21710
rect 49310 21698 49362 21710
rect 6962 21646 6974 21698
rect 7026 21646 7038 21698
rect 7410 21646 7422 21698
rect 7474 21646 7486 21698
rect 7970 21646 7982 21698
rect 8034 21646 8046 21698
rect 11890 21646 11902 21698
rect 11954 21646 11966 21698
rect 19618 21646 19630 21698
rect 19682 21646 19694 21698
rect 23650 21646 23662 21698
rect 23714 21646 23726 21698
rect 26450 21646 26462 21698
rect 26514 21646 26526 21698
rect 28578 21646 28590 21698
rect 28642 21646 28654 21698
rect 31378 21646 31390 21698
rect 31442 21646 31454 21698
rect 36978 21646 36990 21698
rect 37042 21646 37054 21698
rect 45266 21646 45278 21698
rect 45330 21646 45342 21698
rect 47394 21646 47406 21698
rect 47458 21646 47470 21698
rect 14366 21634 14418 21646
rect 24558 21634 24610 21646
rect 42142 21634 42194 21646
rect 49310 21634 49362 21646
rect 51438 21698 51490 21710
rect 56030 21698 56082 21710
rect 53890 21646 53902 21698
rect 53954 21646 53966 21698
rect 54450 21646 54462 21698
rect 54514 21646 54526 21698
rect 57698 21646 57710 21698
rect 57762 21646 57774 21698
rect 51438 21634 51490 21646
rect 56030 21634 56082 21646
rect 3502 21586 3554 21598
rect 13918 21586 13970 21598
rect 16270 21586 16322 21598
rect 1698 21534 1710 21586
rect 1762 21534 1774 21586
rect 3826 21534 3838 21586
rect 3890 21534 3902 21586
rect 6066 21534 6078 21586
rect 6130 21534 6142 21586
rect 7186 21534 7198 21586
rect 7250 21534 7262 21586
rect 8306 21534 8318 21586
rect 8370 21534 8382 21586
rect 8978 21534 8990 21586
rect 9042 21534 9054 21586
rect 10210 21534 10222 21586
rect 10274 21534 10286 21586
rect 10658 21534 10670 21586
rect 10722 21534 10734 21586
rect 11778 21534 11790 21586
rect 11842 21534 11854 21586
rect 16034 21534 16046 21586
rect 16098 21534 16110 21586
rect 3502 21522 3554 21534
rect 13918 21522 13970 21534
rect 16270 21522 16322 21534
rect 17614 21586 17666 21598
rect 20414 21586 20466 21598
rect 23102 21586 23154 21598
rect 25230 21586 25282 21598
rect 31054 21586 31106 21598
rect 38334 21586 38386 21598
rect 42030 21586 42082 21598
rect 17938 21534 17950 21586
rect 18002 21534 18014 21586
rect 19842 21534 19854 21586
rect 19906 21534 19918 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 23874 21534 23886 21586
rect 23938 21534 23950 21586
rect 27682 21534 27694 21586
rect 27746 21534 27758 21586
rect 28690 21534 28702 21586
rect 28754 21534 28766 21586
rect 29698 21534 29710 21586
rect 29762 21534 29774 21586
rect 31826 21534 31838 21586
rect 31890 21534 31902 21586
rect 32274 21534 32286 21586
rect 32338 21534 32350 21586
rect 34402 21534 34414 21586
rect 34466 21534 34478 21586
rect 35858 21534 35870 21586
rect 35922 21534 35934 21586
rect 37538 21534 37550 21586
rect 37602 21534 37614 21586
rect 38770 21534 38782 21586
rect 38834 21534 38846 21586
rect 17614 21522 17666 21534
rect 20414 21522 20466 21534
rect 23102 21522 23154 21534
rect 25230 21522 25282 21534
rect 31054 21522 31106 21534
rect 38334 21522 38386 21534
rect 42030 21522 42082 21534
rect 42366 21586 42418 21598
rect 48750 21586 48802 21598
rect 44034 21534 44046 21586
rect 44098 21534 44110 21586
rect 44706 21534 44718 21586
rect 44770 21534 44782 21586
rect 46610 21534 46622 21586
rect 46674 21534 46686 21586
rect 47170 21534 47182 21586
rect 47234 21534 47246 21586
rect 42366 21522 42418 21534
rect 48750 21522 48802 21534
rect 48974 21586 49026 21598
rect 48974 21522 49026 21534
rect 50990 21586 51042 21598
rect 50990 21522 51042 21534
rect 53342 21586 53394 21598
rect 53342 21522 53394 21534
rect 53790 21586 53842 21598
rect 53790 21522 53842 21534
rect 55246 21586 55298 21598
rect 55246 21522 55298 21534
rect 55470 21586 55522 21598
rect 55794 21534 55806 21586
rect 55858 21534 55870 21586
rect 57250 21534 57262 21586
rect 57314 21534 57326 21586
rect 57922 21534 57934 21586
rect 57986 21534 57998 21586
rect 55470 21522 55522 21534
rect 11454 21474 11506 21486
rect 2706 21422 2718 21474
rect 2770 21422 2782 21474
rect 5954 21422 5966 21474
rect 6018 21422 6030 21474
rect 10322 21422 10334 21474
rect 10386 21422 10398 21474
rect 11454 21410 11506 21422
rect 24334 21474 24386 21486
rect 40238 21474 40290 21486
rect 25666 21422 25678 21474
rect 25730 21422 25742 21474
rect 30146 21422 30158 21474
rect 30210 21422 30222 21474
rect 31938 21422 31950 21474
rect 32002 21422 32014 21474
rect 24334 21410 24386 21422
rect 40238 21410 40290 21422
rect 41134 21474 41186 21486
rect 41134 21410 41186 21422
rect 41470 21474 41522 21486
rect 48190 21474 48242 21486
rect 43698 21422 43710 21474
rect 43762 21422 43774 21474
rect 47618 21422 47630 21474
rect 47682 21422 47694 21474
rect 41470 21410 41522 21422
rect 48190 21410 48242 21422
rect 50654 21474 50706 21486
rect 50654 21410 50706 21422
rect 52782 21474 52834 21486
rect 52782 21410 52834 21422
rect 56702 21474 56754 21486
rect 58034 21422 58046 21474
rect 58098 21422 58110 21474
rect 56702 21410 56754 21422
rect 3390 21362 3442 21374
rect 24670 21362 24722 21374
rect 55694 21362 55746 21374
rect 6402 21310 6414 21362
rect 6466 21310 6478 21362
rect 10098 21310 10110 21362
rect 10162 21310 10174 21362
rect 16034 21310 16046 21362
rect 16098 21310 16110 21362
rect 21410 21310 21422 21362
rect 21474 21310 21486 21362
rect 36754 21310 36766 21362
rect 36818 21310 36830 21362
rect 45042 21310 45054 21362
rect 45106 21310 45118 21362
rect 3390 21298 3442 21310
rect 24670 21298 24722 21310
rect 55694 21298 55746 21310
rect 1344 21194 58576 21228
rect 1344 21142 8367 21194
rect 8419 21142 8471 21194
rect 8523 21142 8575 21194
rect 8627 21142 22674 21194
rect 22726 21142 22778 21194
rect 22830 21142 22882 21194
rect 22934 21142 36981 21194
rect 37033 21142 37085 21194
rect 37137 21142 37189 21194
rect 37241 21142 51288 21194
rect 51340 21142 51392 21194
rect 51444 21142 51496 21194
rect 51548 21142 58576 21194
rect 1344 21108 58576 21142
rect 34862 21026 34914 21038
rect 54350 21026 54402 21038
rect 4946 20974 4958 21026
rect 5010 20974 5022 21026
rect 23650 20974 23662 21026
rect 23714 20974 23726 21026
rect 42130 20974 42142 21026
rect 42194 20974 42206 21026
rect 34862 20962 34914 20974
rect 54350 20962 54402 20974
rect 55246 21026 55298 21038
rect 55246 20962 55298 20974
rect 6302 20914 6354 20926
rect 36430 20914 36482 20926
rect 52894 20914 52946 20926
rect 18498 20862 18510 20914
rect 18562 20862 18574 20914
rect 27010 20862 27022 20914
rect 27074 20862 27086 20914
rect 34514 20862 34526 20914
rect 34578 20862 34590 20914
rect 38546 20862 38558 20914
rect 38610 20862 38622 20914
rect 48066 20862 48078 20914
rect 48130 20862 48142 20914
rect 6302 20850 6354 20862
rect 36430 20850 36482 20862
rect 52894 20850 52946 20862
rect 53790 20914 53842 20926
rect 53790 20850 53842 20862
rect 54798 20914 54850 20926
rect 56466 20862 56478 20914
rect 56530 20862 56542 20914
rect 54798 20850 54850 20862
rect 20414 20802 20466 20814
rect 20750 20802 20802 20814
rect 23998 20802 24050 20814
rect 30382 20802 30434 20814
rect 1810 20750 1822 20802
rect 1874 20750 1886 20802
rect 2594 20750 2606 20802
rect 2658 20750 2670 20802
rect 4722 20750 4734 20802
rect 4786 20750 4798 20802
rect 6738 20750 6750 20802
rect 6802 20750 6814 20802
rect 8418 20750 8430 20802
rect 8482 20750 8494 20802
rect 9650 20750 9662 20802
rect 9714 20750 9726 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 12786 20750 12798 20802
rect 12850 20750 12862 20802
rect 14018 20750 14030 20802
rect 14082 20750 14094 20802
rect 16034 20750 16046 20802
rect 16098 20750 16110 20802
rect 17042 20750 17054 20802
rect 17106 20750 17118 20802
rect 20626 20750 20638 20802
rect 20690 20750 20702 20802
rect 21522 20750 21534 20802
rect 21586 20750 21598 20802
rect 23314 20750 23326 20802
rect 23378 20750 23390 20802
rect 25106 20750 25118 20802
rect 25170 20750 25182 20802
rect 28242 20750 28254 20802
rect 28306 20750 28318 20802
rect 29138 20750 29150 20802
rect 29202 20750 29214 20802
rect 20414 20738 20466 20750
rect 20750 20738 20802 20750
rect 23998 20738 24050 20750
rect 30382 20738 30434 20750
rect 31838 20802 31890 20814
rect 31838 20738 31890 20750
rect 32174 20802 32226 20814
rect 42702 20802 42754 20814
rect 52670 20802 52722 20814
rect 32386 20750 32398 20802
rect 32450 20750 32462 20802
rect 37202 20750 37214 20802
rect 37266 20750 37278 20802
rect 38770 20750 38782 20802
rect 38834 20750 38846 20802
rect 41122 20750 41134 20802
rect 41186 20750 41198 20802
rect 41906 20750 41918 20802
rect 41970 20750 41982 20802
rect 42802 20750 42814 20802
rect 42866 20750 42878 20802
rect 45826 20750 45838 20802
rect 45890 20750 45902 20802
rect 46050 20750 46062 20802
rect 46114 20750 46126 20802
rect 46722 20750 46734 20802
rect 46786 20750 46798 20802
rect 47394 20750 47406 20802
rect 47458 20750 47470 20802
rect 48514 20750 48526 20802
rect 48578 20750 48590 20802
rect 49522 20750 49534 20802
rect 49586 20750 49598 20802
rect 51538 20750 51550 20802
rect 51602 20750 51614 20802
rect 32174 20738 32226 20750
rect 42702 20738 42754 20750
rect 52670 20738 52722 20750
rect 53118 20802 53170 20814
rect 53118 20738 53170 20750
rect 54014 20802 54066 20814
rect 54014 20738 54066 20750
rect 55022 20802 55074 20814
rect 55022 20738 55074 20750
rect 55694 20802 55746 20814
rect 55694 20738 55746 20750
rect 57710 20802 57762 20814
rect 57710 20738 57762 20750
rect 57934 20802 57986 20814
rect 57934 20738 57986 20750
rect 58158 20802 58210 20814
rect 58158 20738 58210 20750
rect 26574 20690 26626 20702
rect 30494 20690 30546 20702
rect 2930 20638 2942 20690
rect 2994 20638 3006 20690
rect 3266 20638 3278 20690
rect 3330 20638 3342 20690
rect 4610 20638 4622 20690
rect 4674 20638 4686 20690
rect 6850 20638 6862 20690
rect 6914 20638 6926 20690
rect 10994 20638 11006 20690
rect 11058 20638 11070 20690
rect 14578 20638 14590 20690
rect 14642 20638 14654 20690
rect 16594 20638 16606 20690
rect 16658 20638 16670 20690
rect 22530 20638 22542 20690
rect 22594 20638 22606 20690
rect 24994 20638 25006 20690
rect 25058 20638 25070 20690
rect 28354 20638 28366 20690
rect 28418 20638 28430 20690
rect 29362 20638 29374 20690
rect 29426 20638 29438 20690
rect 29810 20638 29822 20690
rect 29874 20638 29886 20690
rect 26574 20626 26626 20638
rect 30494 20626 30546 20638
rect 34190 20690 34242 20702
rect 34190 20626 34242 20638
rect 35086 20690 35138 20702
rect 44046 20690 44098 20702
rect 51886 20690 51938 20702
rect 36978 20638 36990 20690
rect 37042 20638 37054 20690
rect 40338 20638 40350 20690
rect 40402 20638 40414 20690
rect 46946 20638 46958 20690
rect 47010 20638 47022 20690
rect 48850 20638 48862 20690
rect 48914 20638 48926 20690
rect 49186 20638 49198 20690
rect 49250 20638 49262 20690
rect 50866 20638 50878 20690
rect 50930 20638 50942 20690
rect 35086 20626 35138 20638
rect 44046 20626 44098 20638
rect 51886 20626 51938 20638
rect 52222 20690 52274 20702
rect 56802 20638 56814 20690
rect 56866 20638 56878 20690
rect 52222 20626 52274 20638
rect 5854 20578 5906 20590
rect 12798 20578 12850 20590
rect 30718 20578 30770 20590
rect 2258 20526 2270 20578
rect 2322 20526 2334 20578
rect 7746 20526 7758 20578
rect 7810 20526 7822 20578
rect 15026 20526 15038 20578
rect 15090 20526 15102 20578
rect 22642 20526 22654 20578
rect 22706 20526 22718 20578
rect 5854 20514 5906 20526
rect 12798 20514 12850 20526
rect 30718 20514 30770 20526
rect 31054 20578 31106 20590
rect 34414 20578 34466 20590
rect 32834 20526 32846 20578
rect 32898 20526 32910 20578
rect 31054 20514 31106 20526
rect 34414 20514 34466 20526
rect 34974 20578 35026 20590
rect 34974 20514 35026 20526
rect 51998 20578 52050 20590
rect 51998 20514 52050 20526
rect 53230 20578 53282 20590
rect 53230 20514 53282 20526
rect 53342 20578 53394 20590
rect 57362 20526 57374 20578
rect 57426 20526 57438 20578
rect 53342 20514 53394 20526
rect 1344 20410 58731 20444
rect 1344 20358 15520 20410
rect 15572 20358 15624 20410
rect 15676 20358 15728 20410
rect 15780 20358 29827 20410
rect 29879 20358 29931 20410
rect 29983 20358 30035 20410
rect 30087 20358 44134 20410
rect 44186 20358 44238 20410
rect 44290 20358 44342 20410
rect 44394 20358 58441 20410
rect 58493 20358 58545 20410
rect 58597 20358 58649 20410
rect 58701 20358 58731 20410
rect 1344 20324 58731 20358
rect 22766 20242 22818 20254
rect 16818 20190 16830 20242
rect 16882 20190 16894 20242
rect 22766 20178 22818 20190
rect 55918 20242 55970 20254
rect 55918 20178 55970 20190
rect 4622 20130 4674 20142
rect 2146 20078 2158 20130
rect 2210 20078 2222 20130
rect 4622 20066 4674 20078
rect 9774 20130 9826 20142
rect 9774 20066 9826 20078
rect 9998 20130 10050 20142
rect 16270 20130 16322 20142
rect 10322 20078 10334 20130
rect 10386 20078 10398 20130
rect 9998 20066 10050 20078
rect 16270 20066 16322 20078
rect 21870 20130 21922 20142
rect 21870 20066 21922 20078
rect 23326 20130 23378 20142
rect 30494 20130 30546 20142
rect 24210 20078 24222 20130
rect 24274 20078 24286 20130
rect 23326 20066 23378 20078
rect 30494 20066 30546 20078
rect 30606 20130 30658 20142
rect 49198 20130 49250 20142
rect 57710 20130 57762 20142
rect 36306 20078 36318 20130
rect 36370 20078 36382 20130
rect 43810 20078 43822 20130
rect 43874 20078 43886 20130
rect 44146 20078 44158 20130
rect 44210 20078 44222 20130
rect 45042 20078 45054 20130
rect 45106 20078 45118 20130
rect 47058 20078 47070 20130
rect 47122 20078 47134 20130
rect 47506 20078 47518 20130
rect 47570 20078 47582 20130
rect 50082 20078 50094 20130
rect 50146 20078 50158 20130
rect 54002 20078 54014 20130
rect 54066 20078 54078 20130
rect 30606 20066 30658 20078
rect 49198 20066 49250 20078
rect 57710 20066 57762 20078
rect 2942 20018 2994 20030
rect 12910 20018 12962 20030
rect 39678 20018 39730 20030
rect 2034 19966 2046 20018
rect 2098 19966 2110 20018
rect 3154 19966 3166 20018
rect 3218 19966 3230 20018
rect 5170 19966 5182 20018
rect 5234 19966 5246 20018
rect 7746 19966 7758 20018
rect 7810 19966 7822 20018
rect 10546 19966 10558 20018
rect 10610 19966 10622 20018
rect 12562 19966 12574 20018
rect 12626 19966 12638 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 15586 19966 15598 20018
rect 15650 19966 15662 20018
rect 17378 19966 17390 20018
rect 17442 19966 17454 20018
rect 21298 19966 21310 20018
rect 21362 19966 21374 20018
rect 24434 19966 24446 20018
rect 24498 19966 24510 20018
rect 25554 19966 25566 20018
rect 25618 19966 25630 20018
rect 25890 19966 25902 20018
rect 25954 19966 25966 20018
rect 27458 19966 27470 20018
rect 27522 19966 27534 20018
rect 28578 19966 28590 20018
rect 28642 19966 28654 20018
rect 30034 19966 30046 20018
rect 30098 19966 30110 20018
rect 33058 19966 33070 20018
rect 33122 19966 33134 20018
rect 34178 19966 34190 20018
rect 34242 19966 34254 20018
rect 35298 19966 35310 20018
rect 35362 19966 35374 20018
rect 36082 19966 36094 20018
rect 36146 19966 36158 20018
rect 37874 19966 37886 20018
rect 37938 19966 37950 20018
rect 2942 19954 2994 19966
rect 12910 19954 12962 19966
rect 39678 19954 39730 19966
rect 40238 20018 40290 20030
rect 47742 20018 47794 20030
rect 42018 19966 42030 20018
rect 42082 19966 42094 20018
rect 42354 19966 42366 20018
rect 42418 19966 42430 20018
rect 44482 19966 44494 20018
rect 44546 19966 44558 20018
rect 46274 19966 46286 20018
rect 46338 19966 46350 20018
rect 40238 19954 40290 19966
rect 47742 19954 47794 19966
rect 49422 20018 49474 20030
rect 55134 20018 55186 20030
rect 50866 19966 50878 20018
rect 50930 19966 50942 20018
rect 51090 19966 51102 20018
rect 51154 19966 51166 20018
rect 52882 19966 52894 20018
rect 52946 19966 52958 20018
rect 53554 19966 53566 20018
rect 53618 19966 53630 20018
rect 53890 19966 53902 20018
rect 53954 19966 53966 20018
rect 49422 19954 49474 19966
rect 55134 19954 55186 19966
rect 55246 20018 55298 20030
rect 55246 19954 55298 19966
rect 55470 20018 55522 20030
rect 55470 19954 55522 19966
rect 56926 20018 56978 20030
rect 56926 19954 56978 19966
rect 7086 19906 7138 19918
rect 9886 19906 9938 19918
rect 16494 19906 16546 19918
rect 21086 19906 21138 19918
rect 38894 19906 38946 19918
rect 4834 19854 4846 19906
rect 4898 19854 4910 19906
rect 7634 19854 7646 19906
rect 7698 19854 7710 19906
rect 8866 19854 8878 19906
rect 8930 19854 8942 19906
rect 15810 19854 15822 19906
rect 15874 19854 15886 19906
rect 19506 19854 19518 19906
rect 19570 19854 19582 19906
rect 37314 19854 37326 19906
rect 37378 19854 37390 19906
rect 7086 19842 7138 19854
rect 9886 19842 9938 19854
rect 16494 19842 16546 19854
rect 21086 19842 21138 19854
rect 38894 19842 38946 19854
rect 39342 19906 39394 19918
rect 43262 19906 43314 19918
rect 41458 19854 41470 19906
rect 41522 19854 41534 19906
rect 39342 19842 39394 19854
rect 43262 19842 43314 19854
rect 48974 19906 49026 19918
rect 48974 19842 49026 19854
rect 49310 19906 49362 19918
rect 49310 19842 49362 19854
rect 2046 19794 2098 19806
rect 23662 19794 23714 19806
rect 30494 19794 30546 19806
rect 48078 19794 48130 19806
rect 10770 19742 10782 19794
rect 10834 19742 10846 19794
rect 29474 19742 29486 19794
rect 29538 19742 29550 19794
rect 35634 19742 35646 19794
rect 35698 19742 35710 19794
rect 46162 19742 46174 19794
rect 46226 19742 46238 19794
rect 2046 19730 2098 19742
rect 23662 19730 23714 19742
rect 30494 19730 30546 19742
rect 48078 19730 48130 19742
rect 48750 19794 48802 19806
rect 48750 19730 48802 19742
rect 1344 19626 58576 19660
rect 1344 19574 8367 19626
rect 8419 19574 8471 19626
rect 8523 19574 8575 19626
rect 8627 19574 22674 19626
rect 22726 19574 22778 19626
rect 22830 19574 22882 19626
rect 22934 19574 36981 19626
rect 37033 19574 37085 19626
rect 37137 19574 37189 19626
rect 37241 19574 51288 19626
rect 51340 19574 51392 19626
rect 51444 19574 51496 19626
rect 51548 19574 58576 19626
rect 1344 19540 58576 19574
rect 11006 19458 11058 19470
rect 23774 19458 23826 19470
rect 15026 19406 15038 19458
rect 15090 19406 15102 19458
rect 11006 19394 11058 19406
rect 23774 19394 23826 19406
rect 26238 19458 26290 19470
rect 36206 19458 36258 19470
rect 45054 19458 45106 19470
rect 35186 19406 35198 19458
rect 35250 19406 35262 19458
rect 43922 19406 43934 19458
rect 43986 19406 43998 19458
rect 45938 19406 45950 19458
rect 46002 19406 46014 19458
rect 53442 19406 53454 19458
rect 53506 19406 53518 19458
rect 26238 19394 26290 19406
rect 36206 19394 36258 19406
rect 45054 19394 45106 19406
rect 19406 19346 19458 19358
rect 15586 19294 15598 19346
rect 15650 19294 15662 19346
rect 16930 19294 16942 19346
rect 16994 19294 17006 19346
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 25106 19294 25118 19346
rect 25170 19294 25182 19346
rect 25890 19294 25902 19346
rect 25954 19294 25966 19346
rect 27010 19294 27022 19346
rect 27074 19294 27086 19346
rect 30258 19294 30270 19346
rect 30322 19294 30334 19346
rect 32386 19294 32398 19346
rect 32450 19294 32462 19346
rect 37538 19294 37550 19346
rect 37602 19294 37614 19346
rect 40562 19294 40574 19346
rect 40626 19294 40638 19346
rect 49634 19294 49646 19346
rect 49698 19294 49710 19346
rect 51650 19294 51662 19346
rect 51714 19294 51726 19346
rect 53106 19294 53118 19346
rect 53170 19294 53182 19346
rect 19406 19282 19458 19294
rect 1710 19234 1762 19246
rect 5742 19234 5794 19246
rect 9326 19234 9378 19246
rect 23326 19234 23378 19246
rect 3602 19182 3614 19234
rect 3666 19182 3678 19234
rect 3938 19182 3950 19234
rect 4002 19182 4014 19234
rect 5842 19182 5854 19234
rect 5906 19182 5918 19234
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 11218 19182 11230 19234
rect 11282 19182 11294 19234
rect 14242 19182 14254 19234
rect 14306 19182 14318 19234
rect 15698 19182 15710 19234
rect 15762 19182 15774 19234
rect 17042 19182 17054 19234
rect 17106 19182 17118 19234
rect 17602 19182 17614 19234
rect 17666 19182 17678 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 1710 19170 1762 19182
rect 5742 19170 5794 19182
rect 9326 19170 9378 19182
rect 23326 19170 23378 19182
rect 23998 19234 24050 19246
rect 29150 19234 29202 19246
rect 35870 19234 35922 19246
rect 47294 19234 47346 19246
rect 53230 19234 53282 19246
rect 24994 19182 25006 19234
rect 25058 19182 25070 19234
rect 25554 19182 25566 19234
rect 25618 19182 25630 19234
rect 27682 19182 27694 19234
rect 27746 19182 27758 19234
rect 29362 19182 29374 19234
rect 29426 19182 29438 19234
rect 31154 19182 31166 19234
rect 31218 19182 31230 19234
rect 32610 19182 32622 19234
rect 32674 19182 32686 19234
rect 33506 19182 33518 19234
rect 33570 19182 33582 19234
rect 34066 19182 34078 19234
rect 34130 19182 34142 19234
rect 37090 19182 37102 19234
rect 37154 19182 37166 19234
rect 38994 19182 39006 19234
rect 39058 19182 39070 19234
rect 41122 19182 41134 19234
rect 41186 19182 41198 19234
rect 41794 19182 41806 19234
rect 41858 19182 41870 19234
rect 43138 19182 43150 19234
rect 43202 19182 43214 19234
rect 46050 19182 46062 19234
rect 46114 19182 46126 19234
rect 47954 19182 47966 19234
rect 48018 19182 48030 19234
rect 49186 19182 49198 19234
rect 49250 19182 49262 19234
rect 49858 19182 49870 19234
rect 49922 19182 49934 19234
rect 50866 19182 50878 19234
rect 50930 19182 50942 19234
rect 53330 19182 53342 19234
rect 53394 19182 53406 19234
rect 54338 19182 54350 19234
rect 54402 19182 54414 19234
rect 58146 19182 58158 19234
rect 58210 19182 58222 19234
rect 23998 19170 24050 19182
rect 29150 19170 29202 19182
rect 35870 19170 35922 19182
rect 47294 19170 47346 19182
rect 53230 19170 53282 19182
rect 2270 19122 2322 19134
rect 7646 19122 7698 19134
rect 16494 19122 16546 19134
rect 4610 19070 4622 19122
rect 4674 19070 4686 19122
rect 8530 19070 8542 19122
rect 8594 19070 8606 19122
rect 8754 19070 8766 19122
rect 8818 19070 8830 19122
rect 10546 19070 10558 19122
rect 10610 19070 10622 19122
rect 11442 19070 11454 19122
rect 11506 19070 11518 19122
rect 2270 19058 2322 19070
rect 7646 19058 7698 19070
rect 16494 19058 16546 19070
rect 18174 19122 18226 19134
rect 18174 19058 18226 19070
rect 23214 19122 23266 19134
rect 26014 19122 26066 19134
rect 36094 19122 36146 19134
rect 45278 19122 45330 19134
rect 57598 19122 57650 19134
rect 24546 19070 24558 19122
rect 24610 19070 24622 19122
rect 28018 19070 28030 19122
rect 28082 19070 28094 19122
rect 33842 19070 33854 19122
rect 33906 19070 33918 19122
rect 37202 19070 37214 19122
rect 37266 19070 37278 19122
rect 40450 19070 40462 19122
rect 40514 19070 40526 19122
rect 43026 19070 43038 19122
rect 43090 19070 43102 19122
rect 49186 19070 49198 19122
rect 49250 19119 49262 19122
rect 49410 19119 49422 19122
rect 49250 19073 49422 19119
rect 49250 19070 49262 19073
rect 49410 19070 49422 19073
rect 49474 19070 49486 19122
rect 54450 19070 54462 19122
rect 54514 19070 54526 19122
rect 56242 19070 56254 19122
rect 56306 19070 56318 19122
rect 23214 19058 23266 19070
rect 26014 19058 26066 19070
rect 36094 19058 36146 19070
rect 45278 19058 45330 19070
rect 57598 19058 57650 19070
rect 5070 19010 5122 19022
rect 20638 19010 20690 19022
rect 9090 18958 9102 19010
rect 9154 18958 9166 19010
rect 19618 18958 19630 19010
rect 19682 18958 19694 19010
rect 5070 18946 5122 18958
rect 20638 18946 20690 18958
rect 22766 19010 22818 19022
rect 22766 18946 22818 18958
rect 24110 19010 24162 19022
rect 24110 18946 24162 18958
rect 45166 19010 45218 19022
rect 49746 18958 49758 19010
rect 49810 18958 49822 19010
rect 45166 18946 45218 18958
rect 1344 18842 58731 18876
rect 1344 18790 15520 18842
rect 15572 18790 15624 18842
rect 15676 18790 15728 18842
rect 15780 18790 29827 18842
rect 29879 18790 29931 18842
rect 29983 18790 30035 18842
rect 30087 18790 44134 18842
rect 44186 18790 44238 18842
rect 44290 18790 44342 18842
rect 44394 18790 58441 18842
rect 58493 18790 58545 18842
rect 58597 18790 58649 18842
rect 58701 18790 58731 18842
rect 1344 18756 58731 18790
rect 2158 18674 2210 18686
rect 2158 18610 2210 18622
rect 4398 18674 4450 18686
rect 26350 18674 26402 18686
rect 14802 18622 14814 18674
rect 14866 18622 14878 18674
rect 4398 18610 4450 18622
rect 26350 18610 26402 18622
rect 26910 18674 26962 18686
rect 35086 18674 35138 18686
rect 28690 18622 28702 18674
rect 28754 18622 28766 18674
rect 26910 18610 26962 18622
rect 35086 18610 35138 18622
rect 35870 18674 35922 18686
rect 35870 18610 35922 18622
rect 39230 18674 39282 18686
rect 39230 18610 39282 18622
rect 41470 18674 41522 18686
rect 41470 18610 41522 18622
rect 41694 18674 41746 18686
rect 45154 18622 45166 18674
rect 45218 18622 45230 18674
rect 51874 18622 51886 18674
rect 51938 18622 51950 18674
rect 41694 18610 41746 18622
rect 19742 18562 19794 18574
rect 26462 18562 26514 18574
rect 34974 18562 35026 18574
rect 3602 18510 3614 18562
rect 3666 18510 3678 18562
rect 3938 18510 3950 18562
rect 4002 18510 4014 18562
rect 5730 18510 5742 18562
rect 5794 18510 5806 18562
rect 6738 18510 6750 18562
rect 6802 18510 6814 18562
rect 14690 18510 14702 18562
rect 14754 18510 14766 18562
rect 18834 18510 18846 18562
rect 18898 18510 18910 18562
rect 23090 18510 23102 18562
rect 23154 18510 23166 18562
rect 25554 18510 25566 18562
rect 25618 18510 25630 18562
rect 28018 18510 28030 18562
rect 28082 18510 28094 18562
rect 19742 18498 19794 18510
rect 26462 18498 26514 18510
rect 34974 18498 35026 18510
rect 35758 18562 35810 18574
rect 41246 18562 41298 18574
rect 37090 18510 37102 18562
rect 37154 18510 37166 18562
rect 44706 18510 44718 18562
rect 44770 18510 44782 18562
rect 48850 18510 48862 18562
rect 48914 18510 48926 18562
rect 52322 18510 52334 18562
rect 52386 18510 52398 18562
rect 54450 18510 54462 18562
rect 54514 18510 54526 18562
rect 35758 18498 35810 18510
rect 41246 18498 41298 18510
rect 2046 18450 2098 18462
rect 4174 18450 4226 18462
rect 2818 18398 2830 18450
rect 2882 18398 2894 18450
rect 3826 18398 3838 18450
rect 3890 18398 3902 18450
rect 2046 18386 2098 18398
rect 4174 18386 4226 18398
rect 4510 18450 4562 18462
rect 4510 18386 4562 18398
rect 5294 18450 5346 18462
rect 8654 18450 8706 18462
rect 26126 18450 26178 18462
rect 6066 18398 6078 18450
rect 6130 18398 6142 18450
rect 6962 18398 6974 18450
rect 7026 18398 7038 18450
rect 9874 18398 9886 18450
rect 9938 18398 9950 18450
rect 10210 18398 10222 18450
rect 10274 18398 10286 18450
rect 11554 18398 11566 18450
rect 11618 18398 11630 18450
rect 11890 18398 11902 18450
rect 11954 18398 11966 18450
rect 13682 18398 13694 18450
rect 13746 18398 13758 18450
rect 15810 18398 15822 18450
rect 15874 18398 15886 18450
rect 17378 18398 17390 18450
rect 17442 18398 17454 18450
rect 18386 18398 18398 18450
rect 18450 18398 18462 18450
rect 20738 18398 20750 18450
rect 20802 18398 20814 18450
rect 22530 18398 22542 18450
rect 22594 18398 22606 18450
rect 25218 18398 25230 18450
rect 25282 18398 25294 18450
rect 5294 18386 5346 18398
rect 8654 18386 8706 18398
rect 26126 18386 26178 18398
rect 27358 18450 27410 18462
rect 29598 18450 29650 18462
rect 33182 18450 33234 18462
rect 29138 18398 29150 18450
rect 29202 18398 29214 18450
rect 30482 18398 30494 18450
rect 30546 18398 30558 18450
rect 30818 18398 30830 18450
rect 30882 18398 30894 18450
rect 27358 18386 27410 18398
rect 29598 18386 29650 18398
rect 33182 18386 33234 18398
rect 33406 18450 33458 18462
rect 33406 18386 33458 18398
rect 33854 18450 33906 18462
rect 33854 18386 33906 18398
rect 36094 18450 36146 18462
rect 36654 18450 36706 18462
rect 42926 18450 42978 18462
rect 54798 18450 54850 18462
rect 36306 18398 36318 18450
rect 36370 18398 36382 18450
rect 37202 18398 37214 18450
rect 37266 18398 37278 18450
rect 38770 18398 38782 18450
rect 38834 18398 38846 18450
rect 42802 18398 42814 18450
rect 42866 18398 42878 18450
rect 43586 18398 43598 18450
rect 43650 18398 43662 18450
rect 45490 18398 45502 18450
rect 45554 18398 45566 18450
rect 46386 18398 46398 18450
rect 46450 18398 46462 18450
rect 46722 18398 46734 18450
rect 46786 18398 46798 18450
rect 47058 18398 47070 18450
rect 47122 18398 47134 18450
rect 49186 18398 49198 18450
rect 49250 18398 49262 18450
rect 50530 18398 50542 18450
rect 50594 18398 50606 18450
rect 52546 18398 52558 18450
rect 52610 18398 52622 18450
rect 53890 18398 53902 18450
rect 53954 18398 53966 18450
rect 36094 18386 36146 18398
rect 36654 18386 36706 18398
rect 42926 18386 42978 18398
rect 54798 18386 54850 18398
rect 54910 18450 54962 18462
rect 54910 18386 54962 18398
rect 2494 18338 2546 18350
rect 11230 18338 11282 18350
rect 20974 18338 21026 18350
rect 6290 18286 6302 18338
rect 6354 18286 6366 18338
rect 8978 18286 8990 18338
rect 9042 18286 9054 18338
rect 9650 18286 9662 18338
rect 9714 18286 9726 18338
rect 18050 18286 18062 18338
rect 18114 18286 18126 18338
rect 2494 18274 2546 18286
rect 11230 18274 11282 18286
rect 20974 18274 21026 18286
rect 21534 18338 21586 18350
rect 34526 18338 34578 18350
rect 22306 18286 22318 18338
rect 22370 18286 22382 18338
rect 24658 18286 24670 18338
rect 24722 18286 24734 18338
rect 25890 18286 25902 18338
rect 25954 18286 25966 18338
rect 30706 18286 30718 18338
rect 30770 18286 30782 18338
rect 21534 18274 21586 18286
rect 34526 18274 34578 18286
rect 36542 18338 36594 18350
rect 36542 18274 36594 18286
rect 40350 18338 40402 18350
rect 40350 18274 40402 18286
rect 41358 18338 41410 18350
rect 41358 18274 41410 18286
rect 42142 18338 42194 18350
rect 55794 18286 55806 18338
rect 55858 18286 55870 18338
rect 42142 18274 42194 18286
rect 16158 18226 16210 18238
rect 33070 18226 33122 18238
rect 7970 18174 7982 18226
rect 8034 18174 8046 18226
rect 10658 18174 10670 18226
rect 10722 18174 10734 18226
rect 22194 18174 22206 18226
rect 22258 18174 22270 18226
rect 31154 18174 31166 18226
rect 31218 18174 31230 18226
rect 16158 18162 16210 18174
rect 33070 18162 33122 18174
rect 33630 18226 33682 18238
rect 33630 18162 33682 18174
rect 35198 18226 35250 18238
rect 35198 18162 35250 18174
rect 42254 18226 42306 18238
rect 42254 18162 42306 18174
rect 1344 18058 58576 18092
rect 1344 18006 8367 18058
rect 8419 18006 8471 18058
rect 8523 18006 8575 18058
rect 8627 18006 22674 18058
rect 22726 18006 22778 18058
rect 22830 18006 22882 18058
rect 22934 18006 36981 18058
rect 37033 18006 37085 18058
rect 37137 18006 37189 18058
rect 37241 18006 51288 18058
rect 51340 18006 51392 18058
rect 51444 18006 51496 18058
rect 51548 18006 58576 18058
rect 1344 17972 58576 18006
rect 28478 17890 28530 17902
rect 42254 17890 42306 17902
rect 19506 17838 19518 17890
rect 19570 17838 19582 17890
rect 32610 17838 32622 17890
rect 32674 17838 32686 17890
rect 28478 17826 28530 17838
rect 42254 17826 42306 17838
rect 43262 17890 43314 17902
rect 43262 17826 43314 17838
rect 2942 17778 2994 17790
rect 4286 17778 4338 17790
rect 7198 17778 7250 17790
rect 3714 17726 3726 17778
rect 3778 17726 3790 17778
rect 6066 17726 6078 17778
rect 6130 17726 6142 17778
rect 2942 17714 2994 17726
rect 4286 17714 4338 17726
rect 7198 17714 7250 17726
rect 11006 17778 11058 17790
rect 11006 17714 11058 17726
rect 12014 17778 12066 17790
rect 40910 17778 40962 17790
rect 45614 17778 45666 17790
rect 15026 17726 15038 17778
rect 15090 17726 15102 17778
rect 17378 17726 17390 17778
rect 17442 17726 17454 17778
rect 20178 17726 20190 17778
rect 20242 17726 20254 17778
rect 39106 17726 39118 17778
rect 39170 17726 39182 17778
rect 41794 17726 41806 17778
rect 41858 17726 41870 17778
rect 42578 17726 42590 17778
rect 42642 17726 42654 17778
rect 45266 17726 45278 17778
rect 45330 17726 45342 17778
rect 12014 17714 12066 17726
rect 40910 17714 40962 17726
rect 45614 17714 45666 17726
rect 53118 17778 53170 17790
rect 53118 17714 53170 17726
rect 57374 17778 57426 17790
rect 57374 17714 57426 17726
rect 2270 17666 2322 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 2270 17602 2322 17614
rect 6862 17666 6914 17678
rect 7982 17666 8034 17678
rect 8318 17666 8370 17678
rect 10446 17666 10498 17678
rect 7074 17614 7086 17666
rect 7138 17614 7150 17666
rect 8194 17614 8206 17666
rect 8258 17614 8270 17666
rect 10210 17614 10222 17666
rect 10274 17614 10286 17666
rect 6862 17602 6914 17614
rect 7982 17602 8034 17614
rect 8318 17602 8370 17614
rect 10446 17602 10498 17614
rect 12350 17666 12402 17678
rect 12350 17602 12402 17614
rect 12910 17666 12962 17678
rect 18174 17666 18226 17678
rect 23774 17666 23826 17678
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 15138 17614 15150 17666
rect 15202 17614 15214 17666
rect 17490 17614 17502 17666
rect 17554 17614 17566 17666
rect 19282 17614 19294 17666
rect 19346 17614 19358 17666
rect 20290 17614 20302 17666
rect 20354 17614 20366 17666
rect 23426 17614 23438 17666
rect 23490 17614 23502 17666
rect 12910 17602 12962 17614
rect 18174 17602 18226 17614
rect 23774 17602 23826 17614
rect 26238 17666 26290 17678
rect 37550 17666 37602 17678
rect 39790 17666 39842 17678
rect 28354 17614 28366 17666
rect 28418 17614 28430 17666
rect 31490 17614 31502 17666
rect 31554 17614 31566 17666
rect 32162 17614 32174 17666
rect 32226 17614 32238 17666
rect 33282 17614 33294 17666
rect 33346 17614 33358 17666
rect 37762 17614 37774 17666
rect 37826 17614 37838 17666
rect 26238 17602 26290 17614
rect 37550 17602 37602 17614
rect 39790 17602 39842 17614
rect 41470 17666 41522 17678
rect 41470 17602 41522 17614
rect 41694 17666 41746 17678
rect 52782 17666 52834 17678
rect 41906 17614 41918 17666
rect 41970 17614 41982 17666
rect 45042 17614 45054 17666
rect 45106 17614 45118 17666
rect 46274 17614 46286 17666
rect 46338 17614 46350 17666
rect 47618 17614 47630 17666
rect 47682 17614 47694 17666
rect 48290 17614 48302 17666
rect 48354 17614 48366 17666
rect 50866 17614 50878 17666
rect 50930 17614 50942 17666
rect 41694 17602 41746 17614
rect 52782 17602 52834 17614
rect 53342 17666 53394 17678
rect 55694 17666 55746 17678
rect 54226 17614 54238 17666
rect 54290 17614 54302 17666
rect 54562 17614 54574 17666
rect 54626 17614 54638 17666
rect 53342 17602 53394 17614
rect 55694 17602 55746 17614
rect 3390 17554 3442 17566
rect 3390 17490 3442 17502
rect 3614 17554 3666 17566
rect 3614 17490 3666 17502
rect 5742 17554 5794 17566
rect 5742 17490 5794 17502
rect 5966 17554 6018 17566
rect 5966 17490 6018 17502
rect 9662 17554 9714 17566
rect 24334 17554 24386 17566
rect 37102 17554 37154 17566
rect 15810 17502 15822 17554
rect 15874 17502 15886 17554
rect 20514 17502 20526 17554
rect 20578 17502 20590 17554
rect 21746 17502 21758 17554
rect 21810 17502 21822 17554
rect 27682 17502 27694 17554
rect 27746 17502 27758 17554
rect 9662 17490 9714 17502
rect 24334 17490 24386 17502
rect 37102 17490 37154 17502
rect 41246 17554 41298 17566
rect 41246 17490 41298 17502
rect 43038 17554 43090 17566
rect 52894 17554 52946 17566
rect 56142 17554 56194 17566
rect 49410 17502 49422 17554
rect 49474 17502 49486 17554
rect 49746 17502 49758 17554
rect 49810 17502 49822 17554
rect 53554 17502 53566 17554
rect 53618 17502 53630 17554
rect 55122 17502 55134 17554
rect 55186 17502 55198 17554
rect 43038 17490 43090 17502
rect 52894 17490 52946 17502
rect 56142 17490 56194 17502
rect 4734 17442 4786 17454
rect 42478 17442 42530 17454
rect 25330 17390 25342 17442
rect 25394 17390 25406 17442
rect 4734 17378 4786 17390
rect 42478 17378 42530 17390
rect 43150 17442 43202 17454
rect 51662 17442 51714 17454
rect 57038 17442 57090 17454
rect 51202 17390 51214 17442
rect 51266 17390 51278 17442
rect 55010 17390 55022 17442
rect 55074 17390 55086 17442
rect 43150 17378 43202 17390
rect 51662 17378 51714 17390
rect 57038 17378 57090 17390
rect 1344 17274 58731 17308
rect 1344 17222 15520 17274
rect 15572 17222 15624 17274
rect 15676 17222 15728 17274
rect 15780 17222 29827 17274
rect 29879 17222 29931 17274
rect 29983 17222 30035 17274
rect 30087 17222 44134 17274
rect 44186 17222 44238 17274
rect 44290 17222 44342 17274
rect 44394 17222 58441 17274
rect 58493 17222 58545 17274
rect 58597 17222 58649 17274
rect 58701 17222 58731 17274
rect 1344 17188 58731 17222
rect 27918 17106 27970 17118
rect 12674 17054 12686 17106
rect 12738 17054 12750 17106
rect 27918 17042 27970 17054
rect 35758 17106 35810 17118
rect 35758 17042 35810 17054
rect 40238 17106 40290 17118
rect 40238 17042 40290 17054
rect 40462 17106 40514 17118
rect 40462 17042 40514 17054
rect 41022 17106 41074 17118
rect 41022 17042 41074 17054
rect 42142 17106 42194 17118
rect 42142 17042 42194 17054
rect 45390 17106 45442 17118
rect 45390 17042 45442 17054
rect 48078 17106 48130 17118
rect 48078 17042 48130 17054
rect 48862 17106 48914 17118
rect 48862 17042 48914 17054
rect 49310 17106 49362 17118
rect 55470 17106 55522 17118
rect 53442 17054 53454 17106
rect 53506 17054 53518 17106
rect 49310 17042 49362 17054
rect 55470 17042 55522 17054
rect 8430 16994 8482 17006
rect 26462 16994 26514 17006
rect 33070 16994 33122 17006
rect 35198 16994 35250 17006
rect 37550 16994 37602 17006
rect 50990 16994 51042 17006
rect 9538 16942 9550 16994
rect 9602 16942 9614 16994
rect 10994 16942 11006 16994
rect 11058 16942 11070 16994
rect 12002 16942 12014 16994
rect 12066 16942 12078 16994
rect 15586 16942 15598 16994
rect 15650 16942 15662 16994
rect 22754 16942 22766 16994
rect 22818 16942 22830 16994
rect 23314 16942 23326 16994
rect 23378 16942 23390 16994
rect 30706 16942 30718 16994
rect 30770 16942 30782 16994
rect 34290 16942 34302 16994
rect 34354 16942 34366 16994
rect 36194 16942 36206 16994
rect 36258 16942 36270 16994
rect 43586 16942 43598 16994
rect 43650 16942 43662 16994
rect 44258 16942 44270 16994
rect 44322 16942 44334 16994
rect 47170 16942 47182 16994
rect 47234 16942 47246 16994
rect 47506 16942 47518 16994
rect 47570 16942 47582 16994
rect 8430 16930 8482 16942
rect 26462 16930 26514 16942
rect 33070 16930 33122 16942
rect 35198 16930 35250 16942
rect 37550 16930 37602 16942
rect 50990 16930 51042 16942
rect 51886 16994 51938 17006
rect 51886 16930 51938 16942
rect 53902 16994 53954 17006
rect 53902 16930 53954 16942
rect 55918 16994 55970 17006
rect 55918 16930 55970 16942
rect 57710 16994 57762 17006
rect 57710 16930 57762 16942
rect 17390 16882 17442 16894
rect 23998 16882 24050 16894
rect 4162 16830 4174 16882
rect 4226 16830 4238 16882
rect 5618 16830 5630 16882
rect 5682 16830 5694 16882
rect 6514 16830 6526 16882
rect 6578 16830 6590 16882
rect 7074 16830 7086 16882
rect 7138 16830 7150 16882
rect 8866 16830 8878 16882
rect 8930 16830 8942 16882
rect 9650 16830 9662 16882
rect 9714 16830 9726 16882
rect 12674 16830 12686 16882
rect 12738 16830 12750 16882
rect 14578 16830 14590 16882
rect 14642 16830 14654 16882
rect 15026 16830 15038 16882
rect 15090 16830 15102 16882
rect 17602 16830 17614 16882
rect 17666 16830 17678 16882
rect 19282 16830 19294 16882
rect 19346 16830 19358 16882
rect 20402 16830 20414 16882
rect 20466 16830 20478 16882
rect 22530 16830 22542 16882
rect 22594 16830 22606 16882
rect 23538 16830 23550 16882
rect 23602 16830 23614 16882
rect 17390 16818 17442 16830
rect 23998 16818 24050 16830
rect 26014 16882 26066 16894
rect 26014 16818 26066 16830
rect 26238 16882 26290 16894
rect 26238 16818 26290 16830
rect 26350 16882 26402 16894
rect 26350 16818 26402 16830
rect 27358 16882 27410 16894
rect 27358 16818 27410 16830
rect 27694 16882 27746 16894
rect 27694 16818 27746 16830
rect 28366 16882 28418 16894
rect 33294 16882 33346 16894
rect 29250 16830 29262 16882
rect 29314 16830 29326 16882
rect 29586 16830 29598 16882
rect 29650 16830 29662 16882
rect 31042 16830 31054 16882
rect 31106 16830 31118 16882
rect 32050 16830 32062 16882
rect 32114 16830 32126 16882
rect 28366 16818 28418 16830
rect 33294 16818 33346 16830
rect 34638 16882 34690 16894
rect 34638 16818 34690 16830
rect 34974 16882 35026 16894
rect 40126 16882 40178 16894
rect 57038 16882 57090 16894
rect 36082 16830 36094 16882
rect 36146 16830 36158 16882
rect 37090 16830 37102 16882
rect 37154 16830 37166 16882
rect 38882 16830 38894 16882
rect 38946 16830 38958 16882
rect 41122 16830 41134 16882
rect 41186 16830 41198 16882
rect 42466 16830 42478 16882
rect 42530 16830 42542 16882
rect 43474 16830 43486 16882
rect 43538 16830 43550 16882
rect 44594 16830 44606 16882
rect 44658 16830 44670 16882
rect 51314 16830 51326 16882
rect 51378 16830 51390 16882
rect 53330 16830 53342 16882
rect 53394 16830 53406 16882
rect 55682 16830 55694 16882
rect 55746 16830 55758 16882
rect 57922 16830 57934 16882
rect 57986 16830 57998 16882
rect 58146 16830 58158 16882
rect 58210 16830 58222 16882
rect 34974 16818 35026 16830
rect 40126 16818 40178 16830
rect 57038 16818 57090 16830
rect 2046 16770 2098 16782
rect 27246 16770 27298 16782
rect 5506 16718 5518 16770
rect 5570 16718 5582 16770
rect 8082 16718 8094 16770
rect 8146 16718 8158 16770
rect 19730 16718 19742 16770
rect 19794 16718 19806 16770
rect 22418 16718 22430 16770
rect 22482 16718 22494 16770
rect 2046 16706 2098 16718
rect 27246 16706 27298 16718
rect 27806 16770 27858 16782
rect 35086 16770 35138 16782
rect 39230 16770 39282 16782
rect 31714 16718 31726 16770
rect 31778 16718 31790 16770
rect 36754 16718 36766 16770
rect 36818 16718 36830 16770
rect 27806 16706 27858 16718
rect 35086 16706 35138 16718
rect 39230 16706 39282 16718
rect 39454 16770 39506 16782
rect 47742 16770 47794 16782
rect 41234 16718 41246 16770
rect 41298 16718 41310 16770
rect 44146 16718 44158 16770
rect 44210 16718 44222 16770
rect 56914 16718 56926 16770
rect 56978 16718 56990 16770
rect 39454 16706 39506 16718
rect 47742 16706 47794 16718
rect 2270 16658 2322 16670
rect 2270 16594 2322 16606
rect 2494 16658 2546 16670
rect 2494 16594 2546 16606
rect 2718 16658 2770 16670
rect 2718 16594 2770 16606
rect 3166 16658 3218 16670
rect 16606 16658 16658 16670
rect 4722 16606 4734 16658
rect 4786 16606 4798 16658
rect 3166 16594 3218 16606
rect 16606 16594 16658 16606
rect 24334 16658 24386 16670
rect 24334 16594 24386 16606
rect 26910 16658 26962 16670
rect 26910 16594 26962 16606
rect 27022 16658 27074 16670
rect 27022 16594 27074 16606
rect 31278 16658 31330 16670
rect 31278 16594 31330 16606
rect 33518 16658 33570 16670
rect 33518 16594 33570 16606
rect 33742 16658 33794 16670
rect 33742 16594 33794 16606
rect 37774 16658 37826 16670
rect 37774 16594 37826 16606
rect 38110 16658 38162 16670
rect 38110 16594 38162 16606
rect 55358 16658 55410 16670
rect 57598 16658 57650 16670
rect 57250 16606 57262 16658
rect 57314 16606 57326 16658
rect 55358 16594 55410 16606
rect 57598 16594 57650 16606
rect 1344 16490 58576 16524
rect 1344 16438 8367 16490
rect 8419 16438 8471 16490
rect 8523 16438 8575 16490
rect 8627 16438 22674 16490
rect 22726 16438 22778 16490
rect 22830 16438 22882 16490
rect 22934 16438 36981 16490
rect 37033 16438 37085 16490
rect 37137 16438 37189 16490
rect 37241 16438 51288 16490
rect 51340 16438 51392 16490
rect 51444 16438 51496 16490
rect 51548 16438 58576 16490
rect 1344 16404 58576 16438
rect 3390 16322 3442 16334
rect 3390 16258 3442 16270
rect 4398 16322 4450 16334
rect 4398 16258 4450 16270
rect 21310 16322 21362 16334
rect 21310 16258 21362 16270
rect 21646 16322 21698 16334
rect 31166 16322 31218 16334
rect 23426 16270 23438 16322
rect 23490 16270 23502 16322
rect 54002 16270 54014 16322
rect 54066 16270 54078 16322
rect 56130 16270 56142 16322
rect 56194 16270 56206 16322
rect 21646 16258 21698 16270
rect 31166 16258 31218 16270
rect 6078 16210 6130 16222
rect 10894 16210 10946 16222
rect 31390 16210 31442 16222
rect 7970 16158 7982 16210
rect 8034 16158 8046 16210
rect 9986 16158 9998 16210
rect 10050 16158 10062 16210
rect 17714 16158 17726 16210
rect 17778 16158 17790 16210
rect 6078 16146 6130 16158
rect 10894 16146 10946 16158
rect 31390 16146 31442 16158
rect 36430 16210 36482 16222
rect 40462 16210 40514 16222
rect 37762 16158 37774 16210
rect 37826 16158 37838 16210
rect 36430 16146 36482 16158
rect 40462 16146 40514 16158
rect 41694 16210 41746 16222
rect 54574 16210 54626 16222
rect 45154 16158 45166 16210
rect 45218 16158 45230 16210
rect 51426 16158 51438 16210
rect 51490 16158 51502 16210
rect 55570 16158 55582 16210
rect 55634 16158 55646 16210
rect 41694 16146 41746 16158
rect 54574 16146 54626 16158
rect 2270 16098 2322 16110
rect 8542 16098 8594 16110
rect 15262 16098 15314 16110
rect 22766 16098 22818 16110
rect 3042 16046 3054 16098
rect 3106 16046 3118 16098
rect 6514 16046 6526 16098
rect 6578 16046 6590 16098
rect 7074 16046 7086 16098
rect 7138 16046 7150 16098
rect 9650 16046 9662 16098
rect 9714 16046 9726 16098
rect 12338 16046 12350 16098
rect 12402 16046 12414 16098
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 17938 16046 17950 16098
rect 18002 16046 18014 16098
rect 18722 16046 18734 16098
rect 18786 16046 18798 16098
rect 20066 16046 20078 16098
rect 20130 16046 20142 16098
rect 22194 16046 22206 16098
rect 22258 16046 22270 16098
rect 2270 16034 2322 16046
rect 8542 16034 8594 16046
rect 15262 16034 15314 16046
rect 22766 16034 22818 16046
rect 23214 16098 23266 16110
rect 26126 16098 26178 16110
rect 24546 16046 24558 16098
rect 24610 16046 24622 16098
rect 23214 16034 23266 16046
rect 26126 16034 26178 16046
rect 26574 16098 26626 16110
rect 30046 16098 30098 16110
rect 27122 16046 27134 16098
rect 27186 16046 27198 16098
rect 27906 16046 27918 16098
rect 27970 16046 27982 16098
rect 28354 16046 28366 16098
rect 28418 16046 28430 16098
rect 26574 16034 26626 16046
rect 30046 16034 30098 16046
rect 30382 16098 30434 16110
rect 38782 16098 38834 16110
rect 36978 16046 36990 16098
rect 37042 16046 37054 16098
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 30382 16034 30434 16046
rect 38782 16034 38834 16046
rect 43710 16098 43762 16110
rect 43710 16034 43762 16046
rect 43934 16098 43986 16110
rect 43934 16034 43986 16046
rect 44382 16098 44434 16110
rect 47854 16098 47906 16110
rect 45042 16046 45054 16098
rect 45106 16046 45118 16098
rect 47618 16046 47630 16098
rect 47682 16046 47694 16098
rect 44382 16034 44434 16046
rect 47854 16034 47906 16046
rect 48974 16098 49026 16110
rect 48974 16034 49026 16046
rect 49310 16098 49362 16110
rect 49310 16034 49362 16046
rect 51102 16098 51154 16110
rect 53678 16098 53730 16110
rect 52098 16046 52110 16098
rect 52162 16046 52174 16098
rect 51102 16034 51154 16046
rect 53678 16034 53730 16046
rect 54910 16098 54962 16110
rect 55794 16046 55806 16098
rect 55858 16046 55870 16098
rect 57362 16046 57374 16098
rect 57426 16046 57438 16098
rect 54910 16034 54962 16046
rect 4622 15986 4674 15998
rect 14478 15986 14530 15998
rect 11218 15934 11230 15986
rect 11282 15934 11294 15986
rect 12674 15934 12686 15986
rect 12738 15934 12750 15986
rect 4622 15922 4674 15934
rect 14478 15922 14530 15934
rect 16606 15986 16658 15998
rect 21534 15986 21586 15998
rect 17154 15934 17166 15986
rect 17218 15934 17230 15986
rect 16606 15922 16658 15934
rect 21534 15922 21586 15934
rect 21982 15986 22034 15998
rect 27358 15986 27410 15998
rect 24322 15934 24334 15986
rect 24386 15934 24398 15986
rect 21982 15922 22034 15934
rect 27358 15922 27410 15934
rect 30158 15986 30210 15998
rect 30158 15922 30210 15934
rect 34862 15986 34914 15998
rect 34862 15922 34914 15934
rect 35086 15986 35138 15998
rect 39230 15986 39282 15998
rect 48078 15986 48130 15998
rect 38210 15934 38222 15986
rect 38274 15934 38286 15986
rect 46498 15934 46510 15986
rect 46562 15934 46574 15986
rect 35086 15922 35138 15934
rect 39230 15922 39282 15934
rect 48078 15922 48130 15934
rect 53230 15986 53282 15998
rect 53230 15922 53282 15934
rect 53454 15986 53506 15998
rect 53454 15922 53506 15934
rect 55022 15986 55074 15998
rect 55022 15922 55074 15934
rect 1710 15874 1762 15886
rect 1710 15810 1762 15822
rect 4510 15874 4562 15886
rect 4510 15810 4562 15822
rect 15038 15874 15090 15886
rect 15038 15810 15090 15822
rect 16270 15874 16322 15886
rect 16270 15810 16322 15822
rect 16494 15874 16546 15886
rect 16494 15810 16546 15822
rect 26686 15874 26738 15886
rect 26686 15810 26738 15822
rect 26910 15874 26962 15886
rect 26910 15810 26962 15822
rect 28478 15874 28530 15886
rect 34974 15874 35026 15886
rect 30818 15822 30830 15874
rect 30882 15822 30894 15874
rect 28478 15810 28530 15822
rect 34974 15810 35026 15822
rect 40238 15874 40290 15886
rect 40238 15810 40290 15822
rect 43822 15874 43874 15886
rect 43822 15810 43874 15822
rect 55246 15874 55298 15886
rect 55246 15810 55298 15822
rect 1344 15706 58731 15740
rect 1344 15654 15520 15706
rect 15572 15654 15624 15706
rect 15676 15654 15728 15706
rect 15780 15654 29827 15706
rect 29879 15654 29931 15706
rect 29983 15654 30035 15706
rect 30087 15654 44134 15706
rect 44186 15654 44238 15706
rect 44290 15654 44342 15706
rect 44394 15654 58441 15706
rect 58493 15654 58545 15706
rect 58597 15654 58649 15706
rect 58701 15654 58731 15706
rect 1344 15620 58731 15654
rect 6750 15538 6802 15550
rect 6750 15474 6802 15486
rect 7422 15538 7474 15550
rect 7422 15474 7474 15486
rect 7870 15538 7922 15550
rect 7870 15474 7922 15486
rect 8878 15538 8930 15550
rect 23102 15538 23154 15550
rect 10098 15486 10110 15538
rect 10162 15486 10174 15538
rect 11554 15486 11566 15538
rect 11618 15486 11630 15538
rect 18722 15486 18734 15538
rect 18786 15486 18798 15538
rect 8878 15474 8930 15486
rect 23102 15474 23154 15486
rect 23326 15538 23378 15550
rect 23326 15474 23378 15486
rect 24446 15538 24498 15550
rect 24446 15474 24498 15486
rect 27918 15538 27970 15550
rect 27918 15474 27970 15486
rect 28142 15538 28194 15550
rect 28142 15474 28194 15486
rect 28254 15538 28306 15550
rect 39006 15538 39058 15550
rect 37090 15486 37102 15538
rect 37154 15486 37166 15538
rect 28254 15474 28306 15486
rect 39006 15474 39058 15486
rect 42142 15538 42194 15550
rect 42142 15474 42194 15486
rect 42590 15538 42642 15550
rect 42590 15474 42642 15486
rect 44606 15538 44658 15550
rect 44606 15474 44658 15486
rect 44830 15538 44882 15550
rect 44830 15474 44882 15486
rect 45390 15538 45442 15550
rect 45390 15474 45442 15486
rect 45838 15538 45890 15550
rect 45838 15474 45890 15486
rect 48078 15538 48130 15550
rect 48078 15474 48130 15486
rect 52110 15538 52162 15550
rect 52110 15474 52162 15486
rect 55246 15538 55298 15550
rect 55246 15474 55298 15486
rect 2606 15426 2658 15438
rect 6638 15426 6690 15438
rect 16046 15426 16098 15438
rect 23886 15426 23938 15438
rect 4386 15374 4398 15426
rect 4450 15374 4462 15426
rect 5282 15374 5294 15426
rect 5346 15374 5358 15426
rect 9650 15374 9662 15426
rect 9714 15374 9726 15426
rect 10546 15374 10558 15426
rect 10610 15374 10622 15426
rect 15474 15374 15486 15426
rect 15538 15374 15550 15426
rect 18050 15374 18062 15426
rect 18114 15374 18126 15426
rect 22306 15374 22318 15426
rect 22370 15374 22382 15426
rect 2606 15362 2658 15374
rect 6638 15362 6690 15374
rect 16046 15362 16098 15374
rect 23886 15362 23938 15374
rect 27022 15426 27074 15438
rect 27022 15362 27074 15374
rect 27694 15426 27746 15438
rect 45726 15426 45778 15438
rect 38098 15374 38110 15426
rect 38162 15374 38174 15426
rect 41682 15374 41694 15426
rect 41746 15374 41758 15426
rect 27694 15362 27746 15374
rect 45726 15362 45778 15374
rect 47854 15426 47906 15438
rect 47854 15362 47906 15374
rect 50654 15426 50706 15438
rect 50654 15362 50706 15374
rect 50990 15426 51042 15438
rect 54674 15374 54686 15426
rect 54738 15374 54750 15426
rect 58034 15374 58046 15426
rect 58098 15374 58110 15426
rect 50990 15362 51042 15374
rect 2382 15314 2434 15326
rect 2382 15250 2434 15262
rect 3054 15314 3106 15326
rect 6974 15314 7026 15326
rect 16270 15314 16322 15326
rect 6066 15262 6078 15314
rect 6130 15262 6142 15314
rect 8978 15262 8990 15314
rect 9042 15262 9054 15314
rect 9538 15262 9550 15314
rect 9602 15262 9614 15314
rect 10658 15262 10670 15314
rect 10722 15262 10734 15314
rect 11442 15262 11454 15314
rect 11506 15262 11518 15314
rect 12338 15262 12350 15314
rect 12402 15262 12414 15314
rect 13906 15262 13918 15314
rect 13970 15262 13982 15314
rect 14130 15262 14142 15314
rect 14194 15262 14206 15314
rect 3054 15250 3106 15262
rect 6974 15250 7026 15262
rect 16270 15250 16322 15262
rect 16382 15314 16434 15326
rect 23438 15314 23490 15326
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 18610 15262 18622 15314
rect 18674 15262 18686 15314
rect 19170 15262 19182 15314
rect 19234 15262 19246 15314
rect 19506 15262 19518 15314
rect 19570 15262 19582 15314
rect 21522 15262 21534 15314
rect 21586 15262 21598 15314
rect 16382 15250 16434 15262
rect 23438 15250 23490 15262
rect 25230 15314 25282 15326
rect 30830 15314 30882 15326
rect 32510 15314 32562 15326
rect 25442 15262 25454 15314
rect 25506 15262 25518 15314
rect 31042 15262 31054 15314
rect 31106 15262 31118 15314
rect 32050 15262 32062 15314
rect 32114 15262 32126 15314
rect 25230 15250 25282 15262
rect 30830 15250 30882 15262
rect 32510 15250 32562 15262
rect 33966 15314 34018 15326
rect 33966 15250 34018 15262
rect 34190 15314 34242 15326
rect 34190 15250 34242 15262
rect 34414 15314 34466 15326
rect 34414 15250 34466 15262
rect 34638 15314 34690 15326
rect 34638 15250 34690 15262
rect 34974 15314 35026 15326
rect 42366 15314 42418 15326
rect 35186 15262 35198 15314
rect 35250 15262 35262 15314
rect 36978 15262 36990 15314
rect 37042 15262 37054 15314
rect 37874 15262 37886 15314
rect 37938 15262 37950 15314
rect 41122 15262 41134 15314
rect 41186 15262 41198 15314
rect 34974 15250 35026 15262
rect 42366 15250 42418 15262
rect 44270 15314 44322 15326
rect 44270 15250 44322 15262
rect 47518 15314 47570 15326
rect 51214 15314 51266 15326
rect 48962 15262 48974 15314
rect 49026 15262 49038 15314
rect 49186 15262 49198 15314
rect 49250 15262 49262 15314
rect 47518 15250 47570 15262
rect 51214 15250 51266 15262
rect 51438 15314 51490 15326
rect 51438 15250 51490 15262
rect 51662 15314 51714 15326
rect 51662 15250 51714 15262
rect 53454 15314 53506 15326
rect 53454 15250 53506 15262
rect 53678 15314 53730 15326
rect 53678 15250 53730 15262
rect 54126 15314 54178 15326
rect 57138 15262 57150 15314
rect 57202 15262 57214 15314
rect 54126 15250 54178 15262
rect 24110 15202 24162 15214
rect 33518 15202 33570 15214
rect 39342 15202 39394 15214
rect 42478 15202 42530 15214
rect 48750 15202 48802 15214
rect 2034 15150 2046 15202
rect 2098 15150 2110 15202
rect 14242 15150 14254 15202
rect 14306 15150 14318 15202
rect 22082 15150 22094 15202
rect 22146 15150 22158 15202
rect 28242 15150 28254 15202
rect 28306 15150 28318 15202
rect 31714 15150 31726 15202
rect 31778 15150 31790 15202
rect 38322 15150 38334 15202
rect 38386 15150 38398 15202
rect 41570 15150 41582 15202
rect 41634 15150 41646 15202
rect 48178 15150 48190 15202
rect 48242 15150 48254 15202
rect 24110 15138 24162 15150
rect 33518 15138 33570 15150
rect 39342 15138 39394 15150
rect 42478 15138 42530 15150
rect 48750 15138 48802 15150
rect 53902 15202 53954 15214
rect 53902 15138 53954 15150
rect 55806 15202 55858 15214
rect 55806 15138 55858 15150
rect 6078 15090 6130 15102
rect 44494 15090 44546 15102
rect 7074 15038 7086 15090
rect 7138 15087 7150 15090
rect 7410 15087 7422 15090
rect 7138 15041 7422 15087
rect 7138 15038 7150 15041
rect 7410 15038 7422 15041
rect 7474 15038 7486 15090
rect 7634 15038 7646 15090
rect 7698 15087 7710 15090
rect 7970 15087 7982 15090
rect 7698 15041 7982 15087
rect 7698 15038 7710 15041
rect 7970 15038 7982 15041
rect 8034 15038 8046 15090
rect 35634 15038 35646 15090
rect 35698 15038 35710 15090
rect 6078 15026 6130 15038
rect 44494 15026 44546 15038
rect 45838 15090 45890 15102
rect 45838 15026 45890 15038
rect 1344 14922 58576 14956
rect 1344 14870 8367 14922
rect 8419 14870 8471 14922
rect 8523 14870 8575 14922
rect 8627 14870 22674 14922
rect 22726 14870 22778 14922
rect 22830 14870 22882 14922
rect 22934 14870 36981 14922
rect 37033 14870 37085 14922
rect 37137 14870 37189 14922
rect 37241 14870 51288 14922
rect 51340 14870 51392 14922
rect 51444 14870 51496 14922
rect 51548 14870 58576 14922
rect 1344 14836 58576 14870
rect 8654 14754 8706 14766
rect 24222 14754 24274 14766
rect 8978 14702 8990 14754
rect 9042 14702 9054 14754
rect 8654 14690 8706 14702
rect 24222 14690 24274 14702
rect 28366 14754 28418 14766
rect 33506 14702 33518 14754
rect 33570 14702 33582 14754
rect 38658 14702 38670 14754
rect 38722 14702 38734 14754
rect 28366 14690 28418 14702
rect 6302 14642 6354 14654
rect 8430 14642 8482 14654
rect 13582 14642 13634 14654
rect 23662 14642 23714 14654
rect 7634 14590 7646 14642
rect 7698 14590 7710 14642
rect 12114 14590 12126 14642
rect 12178 14590 12190 14642
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 21858 14590 21870 14642
rect 21922 14590 21934 14642
rect 22418 14590 22430 14642
rect 22482 14590 22494 14642
rect 6302 14578 6354 14590
rect 8430 14578 8482 14590
rect 13582 14578 13634 14590
rect 23662 14578 23714 14590
rect 23886 14642 23938 14654
rect 53454 14642 53506 14654
rect 33058 14590 33070 14642
rect 33122 14590 33134 14642
rect 34738 14590 34750 14642
rect 34802 14590 34814 14642
rect 37874 14590 37886 14642
rect 37938 14590 37950 14642
rect 39554 14590 39566 14642
rect 39618 14590 39630 14642
rect 41458 14590 41470 14642
rect 41522 14590 41534 14642
rect 23886 14578 23938 14590
rect 53454 14578 53506 14590
rect 2606 14530 2658 14542
rect 2606 14466 2658 14478
rect 2942 14530 2994 14542
rect 4286 14530 4338 14542
rect 10782 14530 10834 14542
rect 3938 14478 3950 14530
rect 4002 14478 4014 14530
rect 7522 14478 7534 14530
rect 7586 14478 7598 14530
rect 2942 14466 2994 14478
rect 4286 14466 4338 14478
rect 10782 14466 10834 14478
rect 11006 14530 11058 14542
rect 11006 14466 11058 14478
rect 11342 14530 11394 14542
rect 22878 14530 22930 14542
rect 11554 14478 11566 14530
rect 11618 14478 11630 14530
rect 12226 14478 12238 14530
rect 12290 14478 12302 14530
rect 16034 14478 16046 14530
rect 16098 14478 16110 14530
rect 18162 14478 18174 14530
rect 18226 14478 18238 14530
rect 18610 14478 18622 14530
rect 18674 14478 18686 14530
rect 21634 14478 21646 14530
rect 21698 14478 21710 14530
rect 22642 14478 22654 14530
rect 22706 14478 22718 14530
rect 11342 14466 11394 14478
rect 22878 14466 22930 14478
rect 24446 14530 24498 14542
rect 27470 14530 27522 14542
rect 24770 14478 24782 14530
rect 24834 14478 24846 14530
rect 24446 14466 24498 14478
rect 27470 14466 27522 14478
rect 30718 14530 30770 14542
rect 35758 14530 35810 14542
rect 40574 14530 40626 14542
rect 31154 14478 31166 14530
rect 31218 14478 31230 14530
rect 32946 14478 32958 14530
rect 33010 14478 33022 14530
rect 34850 14478 34862 14530
rect 34914 14478 34926 14530
rect 37986 14478 37998 14530
rect 38050 14478 38062 14530
rect 38210 14478 38222 14530
rect 38274 14478 38286 14530
rect 30718 14466 30770 14478
rect 35758 14466 35810 14478
rect 40574 14466 40626 14478
rect 41358 14530 41410 14542
rect 44830 14530 44882 14542
rect 41682 14478 41694 14530
rect 41746 14478 41758 14530
rect 41358 14466 41410 14478
rect 44830 14466 44882 14478
rect 45054 14530 45106 14542
rect 50878 14530 50930 14542
rect 48178 14478 48190 14530
rect 48242 14478 48254 14530
rect 49186 14478 49198 14530
rect 49250 14478 49262 14530
rect 45054 14466 45106 14478
rect 50878 14466 50930 14478
rect 51214 14530 51266 14542
rect 51214 14466 51266 14478
rect 51438 14530 51490 14542
rect 51438 14466 51490 14478
rect 53006 14530 53058 14542
rect 53006 14466 53058 14478
rect 53230 14530 53282 14542
rect 53230 14466 53282 14478
rect 54462 14530 54514 14542
rect 54462 14466 54514 14478
rect 56478 14530 56530 14542
rect 56478 14466 56530 14478
rect 2270 14418 2322 14430
rect 2270 14354 2322 14366
rect 4398 14418 4450 14430
rect 4398 14354 4450 14366
rect 4734 14418 4786 14430
rect 4734 14354 4786 14366
rect 8094 14418 8146 14430
rect 8094 14354 8146 14366
rect 9550 14418 9602 14430
rect 14254 14418 14306 14430
rect 16382 14418 16434 14430
rect 12898 14366 12910 14418
rect 12962 14366 12974 14418
rect 14578 14366 14590 14418
rect 14642 14366 14654 14418
rect 9550 14354 9602 14366
rect 14254 14354 14306 14366
rect 16382 14354 16434 14366
rect 17166 14418 17218 14430
rect 17166 14354 17218 14366
rect 19742 14418 19794 14430
rect 19742 14354 19794 14366
rect 23214 14418 23266 14430
rect 27134 14418 27186 14430
rect 26002 14366 26014 14418
rect 26066 14366 26078 14418
rect 23214 14354 23266 14366
rect 27134 14354 27186 14366
rect 28366 14418 28418 14430
rect 28366 14354 28418 14366
rect 28478 14418 28530 14430
rect 28478 14354 28530 14366
rect 35870 14418 35922 14430
rect 35870 14354 35922 14366
rect 39230 14418 39282 14430
rect 39230 14354 39282 14366
rect 45278 14418 45330 14430
rect 55022 14418 55074 14430
rect 47506 14366 47518 14418
rect 47570 14366 47582 14418
rect 49074 14366 49086 14418
rect 49138 14366 49150 14418
rect 45278 14354 45330 14366
rect 55022 14354 55074 14366
rect 57038 14418 57090 14430
rect 57038 14354 57090 14366
rect 1710 14306 1762 14318
rect 1710 14242 1762 14254
rect 2718 14306 2770 14318
rect 2718 14242 2770 14254
rect 4846 14306 4898 14318
rect 4846 14242 4898 14254
rect 5070 14306 5122 14318
rect 5070 14242 5122 14254
rect 5854 14306 5906 14318
rect 5854 14242 5906 14254
rect 9214 14306 9266 14318
rect 9214 14242 9266 14254
rect 9438 14306 9490 14318
rect 9438 14242 9490 14254
rect 10446 14306 10498 14318
rect 10446 14242 10498 14254
rect 11118 14306 11170 14318
rect 11118 14242 11170 14254
rect 23102 14306 23154 14318
rect 23102 14242 23154 14254
rect 26798 14306 26850 14318
rect 26798 14242 26850 14254
rect 27246 14306 27298 14318
rect 27246 14242 27298 14254
rect 27806 14306 27858 14318
rect 27806 14242 27858 14254
rect 34750 14306 34802 14318
rect 34750 14242 34802 14254
rect 36094 14306 36146 14318
rect 36094 14242 36146 14254
rect 39454 14306 39506 14318
rect 39454 14242 39506 14254
rect 40686 14306 40738 14318
rect 40686 14242 40738 14254
rect 40910 14306 40962 14318
rect 44942 14306 44994 14318
rect 49982 14306 50034 14318
rect 41906 14254 41918 14306
rect 41970 14254 41982 14306
rect 48514 14254 48526 14306
rect 48578 14254 48590 14306
rect 40910 14242 40962 14254
rect 44942 14242 44994 14254
rect 49982 14242 50034 14254
rect 50542 14306 50594 14318
rect 50542 14242 50594 14254
rect 51102 14306 51154 14318
rect 51102 14242 51154 14254
rect 52110 14306 52162 14318
rect 52110 14242 52162 14254
rect 52558 14306 52610 14318
rect 54562 14254 54574 14306
rect 54626 14254 54638 14306
rect 52558 14242 52610 14254
rect 1344 14138 58731 14172
rect 1344 14086 15520 14138
rect 15572 14086 15624 14138
rect 15676 14086 15728 14138
rect 15780 14086 29827 14138
rect 29879 14086 29931 14138
rect 29983 14086 30035 14138
rect 30087 14086 44134 14138
rect 44186 14086 44238 14138
rect 44290 14086 44342 14138
rect 44394 14086 58441 14138
rect 58493 14086 58545 14138
rect 58597 14086 58649 14138
rect 58701 14086 58731 14138
rect 1344 14052 58731 14086
rect 6638 13970 6690 13982
rect 5730 13918 5742 13970
rect 5794 13918 5806 13970
rect 6638 13906 6690 13918
rect 6750 13970 6802 13982
rect 6750 13906 6802 13918
rect 6862 13970 6914 13982
rect 6862 13906 6914 13918
rect 9550 13970 9602 13982
rect 9550 13906 9602 13918
rect 13806 13970 13858 13982
rect 13806 13906 13858 13918
rect 15710 13970 15762 13982
rect 15710 13906 15762 13918
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 18174 13970 18226 13982
rect 23326 13970 23378 13982
rect 22530 13918 22542 13970
rect 22594 13918 22606 13970
rect 18174 13906 18226 13918
rect 23326 13906 23378 13918
rect 23774 13970 23826 13982
rect 23774 13906 23826 13918
rect 25902 13970 25954 13982
rect 25902 13906 25954 13918
rect 26798 13970 26850 13982
rect 26798 13906 26850 13918
rect 27694 13970 27746 13982
rect 27694 13906 27746 13918
rect 28478 13970 28530 13982
rect 28478 13906 28530 13918
rect 29262 13970 29314 13982
rect 45054 13970 45106 13982
rect 51214 13970 51266 13982
rect 30706 13918 30718 13970
rect 30770 13918 30782 13970
rect 34402 13918 34414 13970
rect 34466 13918 34478 13970
rect 49298 13918 49310 13970
rect 49362 13918 49374 13970
rect 29262 13906 29314 13918
rect 45054 13906 45106 13918
rect 51214 13906 51266 13918
rect 55806 13970 55858 13982
rect 55806 13906 55858 13918
rect 55918 13970 55970 13982
rect 55918 13906 55970 13918
rect 2830 13858 2882 13870
rect 12350 13858 12402 13870
rect 16718 13858 16770 13870
rect 5954 13806 5966 13858
rect 6018 13806 6030 13858
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 15026 13806 15038 13858
rect 15090 13806 15102 13858
rect 2830 13794 2882 13806
rect 12350 13794 12402 13806
rect 16718 13794 16770 13806
rect 21982 13858 22034 13870
rect 21982 13794 22034 13806
rect 28702 13858 28754 13870
rect 28702 13794 28754 13806
rect 28814 13858 28866 13870
rect 36094 13858 36146 13870
rect 30034 13806 30046 13858
rect 30098 13806 30110 13858
rect 28814 13794 28866 13806
rect 36094 13794 36146 13806
rect 41582 13858 41634 13870
rect 41582 13794 41634 13806
rect 44606 13858 44658 13870
rect 44606 13794 44658 13806
rect 45502 13858 45554 13870
rect 51662 13858 51714 13870
rect 48850 13806 48862 13858
rect 48914 13806 48926 13858
rect 50306 13806 50318 13858
rect 50370 13806 50382 13858
rect 45502 13794 45554 13806
rect 51662 13794 51714 13806
rect 4286 13746 4338 13758
rect 3938 13694 3950 13746
rect 4002 13694 4014 13746
rect 4286 13682 4338 13694
rect 6190 13746 6242 13758
rect 10446 13746 10498 13758
rect 7634 13694 7646 13746
rect 7698 13694 7710 13746
rect 7858 13694 7870 13746
rect 7922 13694 7934 13746
rect 8978 13694 8990 13746
rect 9042 13694 9054 13746
rect 6190 13682 6242 13694
rect 10446 13682 10498 13694
rect 11118 13746 11170 13758
rect 16158 13746 16210 13758
rect 25342 13746 25394 13758
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 11666 13694 11678 13746
rect 11730 13694 11742 13746
rect 12674 13694 12686 13746
rect 12738 13694 12750 13746
rect 17602 13694 17614 13746
rect 17666 13694 17678 13746
rect 18946 13694 18958 13746
rect 19010 13694 19022 13746
rect 21186 13694 21198 13746
rect 21250 13694 21262 13746
rect 11118 13682 11170 13694
rect 16158 13682 16210 13694
rect 25342 13682 25394 13694
rect 26686 13746 26738 13758
rect 26686 13682 26738 13694
rect 26910 13746 26962 13758
rect 26910 13682 26962 13694
rect 27806 13746 27858 13758
rect 27806 13682 27858 13694
rect 27918 13746 27970 13758
rect 27918 13682 27970 13694
rect 28366 13746 28418 13758
rect 35758 13746 35810 13758
rect 41358 13746 41410 13758
rect 30258 13694 30270 13746
rect 30322 13694 30334 13746
rect 36754 13694 36766 13746
rect 36818 13694 36830 13746
rect 37426 13694 37438 13746
rect 37490 13694 37502 13746
rect 40114 13694 40126 13746
rect 40178 13694 40190 13746
rect 28366 13682 28418 13694
rect 35758 13682 35810 13694
rect 41358 13682 41410 13694
rect 42030 13746 42082 13758
rect 44830 13746 44882 13758
rect 49870 13746 49922 13758
rect 42242 13694 42254 13746
rect 42306 13694 42318 13746
rect 45714 13694 45726 13746
rect 45778 13694 45790 13746
rect 48738 13694 48750 13746
rect 48802 13694 48814 13746
rect 42030 13682 42082 13694
rect 44830 13682 44882 13694
rect 49870 13682 49922 13694
rect 52558 13746 52610 13758
rect 52558 13682 52610 13694
rect 54350 13746 54402 13758
rect 54350 13682 54402 13694
rect 54798 13746 54850 13758
rect 54798 13682 54850 13694
rect 55358 13746 55410 13758
rect 55358 13682 55410 13694
rect 56030 13746 56082 13758
rect 57586 13694 57598 13746
rect 57650 13694 57662 13746
rect 56030 13682 56082 13694
rect 1934 13634 1986 13646
rect 1934 13570 1986 13582
rect 9662 13634 9714 13646
rect 9662 13570 9714 13582
rect 10670 13634 10722 13646
rect 18622 13634 18674 13646
rect 24334 13634 24386 13646
rect 12786 13582 12798 13634
rect 12850 13582 12862 13634
rect 18946 13631 18958 13634
rect 10670 13570 10722 13582
rect 18622 13570 18674 13582
rect 18737 13585 18958 13631
rect 8766 13522 8818 13534
rect 8766 13458 8818 13470
rect 10334 13522 10386 13534
rect 10334 13458 10386 13470
rect 10782 13522 10834 13534
rect 10782 13458 10834 13470
rect 15374 13522 15426 13534
rect 18737 13522 18783 13585
rect 18946 13582 18958 13585
rect 19010 13582 19022 13634
rect 21074 13582 21086 13634
rect 21138 13582 21150 13634
rect 24334 13570 24386 13582
rect 24670 13634 24722 13646
rect 24670 13570 24722 13582
rect 25230 13634 25282 13646
rect 25230 13570 25282 13582
rect 26462 13634 26514 13646
rect 26462 13570 26514 13582
rect 29710 13634 29762 13646
rect 29710 13570 29762 13582
rect 34750 13634 34802 13646
rect 34750 13570 34802 13582
rect 34974 13634 35026 13646
rect 34974 13570 35026 13582
rect 35870 13634 35922 13646
rect 42926 13634 42978 13646
rect 37874 13582 37886 13634
rect 37938 13582 37950 13634
rect 39554 13582 39566 13634
rect 39618 13582 39630 13634
rect 35870 13570 35922 13582
rect 42926 13570 42978 13582
rect 44158 13634 44210 13646
rect 44158 13570 44210 13582
rect 44942 13634 44994 13646
rect 44942 13570 44994 13582
rect 52894 13634 52946 13646
rect 58158 13634 58210 13646
rect 57250 13582 57262 13634
rect 57314 13582 57326 13634
rect 52894 13570 52946 13582
rect 58158 13570 58210 13582
rect 22206 13522 22258 13534
rect 18722 13470 18734 13522
rect 18786 13470 18798 13522
rect 21522 13470 21534 13522
rect 21586 13470 21598 13522
rect 15374 13458 15426 13470
rect 22206 13458 22258 13470
rect 26238 13522 26290 13534
rect 26238 13458 26290 13470
rect 41022 13522 41074 13534
rect 41022 13458 41074 13470
rect 45390 13522 45442 13534
rect 55010 13470 55022 13522
rect 55074 13470 55086 13522
rect 45390 13458 45442 13470
rect 1344 13354 58576 13388
rect 1344 13302 8367 13354
rect 8419 13302 8471 13354
rect 8523 13302 8575 13354
rect 8627 13302 22674 13354
rect 22726 13302 22778 13354
rect 22830 13302 22882 13354
rect 22934 13302 36981 13354
rect 37033 13302 37085 13354
rect 37137 13302 37189 13354
rect 37241 13302 51288 13354
rect 51340 13302 51392 13354
rect 51444 13302 51496 13354
rect 51548 13302 58576 13354
rect 1344 13268 58576 13302
rect 2718 13186 2770 13198
rect 17950 13186 18002 13198
rect 12226 13134 12238 13186
rect 12290 13134 12302 13186
rect 2718 13122 2770 13134
rect 17950 13122 18002 13134
rect 19630 13186 19682 13198
rect 30942 13186 30994 13198
rect 28242 13134 28254 13186
rect 28306 13134 28318 13186
rect 19630 13122 19682 13134
rect 30942 13122 30994 13134
rect 46174 13186 46226 13198
rect 46174 13122 46226 13134
rect 47294 13186 47346 13198
rect 47294 13122 47346 13134
rect 48750 13186 48802 13198
rect 48750 13122 48802 13134
rect 49086 13186 49138 13198
rect 53118 13186 53170 13198
rect 49970 13134 49982 13186
rect 50034 13183 50046 13186
rect 50034 13137 50815 13183
rect 50034 13134 50046 13137
rect 49086 13122 49138 13134
rect 5966 13074 6018 13086
rect 9886 13074 9938 13086
rect 4386 13022 4398 13074
rect 4450 13022 4462 13074
rect 4834 13022 4846 13074
rect 4898 13022 4910 13074
rect 8306 13022 8318 13074
rect 8370 13022 8382 13074
rect 5966 13010 6018 13022
rect 9886 13010 9938 13022
rect 10334 13074 10386 13086
rect 10334 13010 10386 13022
rect 11118 13074 11170 13086
rect 11118 13010 11170 13022
rect 14254 13074 14306 13086
rect 14254 13010 14306 13022
rect 15374 13074 15426 13086
rect 15374 13010 15426 13022
rect 16270 13074 16322 13086
rect 16270 13010 16322 13022
rect 19294 13074 19346 13086
rect 19294 13010 19346 13022
rect 20638 13074 20690 13086
rect 22990 13074 23042 13086
rect 45166 13074 45218 13086
rect 21410 13022 21422 13074
rect 21474 13022 21486 13074
rect 24770 13022 24782 13074
rect 24834 13022 24846 13074
rect 28354 13022 28366 13074
rect 28418 13022 28430 13074
rect 20638 13010 20690 13022
rect 22990 13010 23042 13022
rect 45166 13010 45218 13022
rect 46734 13074 46786 13086
rect 50318 13074 50370 13086
rect 47618 13022 47630 13074
rect 47682 13022 47694 13074
rect 46734 13010 46786 13022
rect 50318 13010 50370 13022
rect 11006 12962 11058 12974
rect 1922 12910 1934 12962
rect 1986 12910 1998 12962
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 5058 12910 5070 12962
rect 5122 12910 5134 12962
rect 8194 12910 8206 12962
rect 8258 12910 8270 12962
rect 11006 12898 11058 12910
rect 11342 12962 11394 12974
rect 14814 12962 14866 12974
rect 11666 12910 11678 12962
rect 11730 12910 11742 12962
rect 12226 12910 12238 12962
rect 12290 12910 12302 12962
rect 12562 12910 12574 12962
rect 12626 12910 12638 12962
rect 11342 12898 11394 12910
rect 14814 12898 14866 12910
rect 17614 12962 17666 12974
rect 20190 12962 20242 12974
rect 26910 12962 26962 12974
rect 35310 12962 35362 12974
rect 18610 12910 18622 12962
rect 18674 12910 18686 12962
rect 21858 12910 21870 12962
rect 21922 12910 21934 12962
rect 23314 12910 23326 12962
rect 23378 12910 23390 12962
rect 27234 12910 27246 12962
rect 27298 12910 27310 12962
rect 28130 12910 28142 12962
rect 28194 12910 28206 12962
rect 30594 12910 30606 12962
rect 30658 12910 30670 12962
rect 31266 12910 31278 12962
rect 31330 12910 31342 12962
rect 33282 12910 33294 12962
rect 33346 12910 33358 12962
rect 17614 12898 17666 12910
rect 20190 12898 20242 12910
rect 26910 12898 26962 12910
rect 35310 12898 35362 12910
rect 35870 12962 35922 12974
rect 37774 12962 37826 12974
rect 45502 12962 45554 12974
rect 37314 12910 37326 12962
rect 37378 12959 37390 12962
rect 37538 12959 37550 12962
rect 37378 12913 37550 12959
rect 37378 12910 37390 12913
rect 37538 12910 37550 12913
rect 37602 12910 37614 12962
rect 38546 12910 38558 12962
rect 38610 12910 38622 12962
rect 39890 12910 39902 12962
rect 39954 12910 39966 12962
rect 40338 12910 40350 12962
rect 40402 12910 40414 12962
rect 35870 12898 35922 12910
rect 37774 12898 37826 12910
rect 45502 12898 45554 12910
rect 48078 12962 48130 12974
rect 48078 12898 48130 12910
rect 48526 12962 48578 12974
rect 48526 12898 48578 12910
rect 48974 12962 49026 12974
rect 48974 12898 49026 12910
rect 10670 12850 10722 12862
rect 9426 12798 9438 12850
rect 9490 12798 9502 12850
rect 10670 12786 10722 12798
rect 15486 12850 15538 12862
rect 15486 12786 15538 12798
rect 15934 12850 15986 12862
rect 15934 12786 15986 12798
rect 16382 12850 16434 12862
rect 22318 12850 22370 12862
rect 33854 12850 33906 12862
rect 17042 12798 17054 12850
rect 17106 12798 17118 12850
rect 17378 12798 17390 12850
rect 17442 12798 17454 12850
rect 18498 12798 18510 12850
rect 18562 12798 18574 12850
rect 31378 12798 31390 12850
rect 31442 12798 31454 12850
rect 16382 12786 16434 12798
rect 22318 12786 22370 12798
rect 33854 12786 33906 12798
rect 35758 12850 35810 12862
rect 35758 12786 35810 12798
rect 37662 12850 37714 12862
rect 41234 12798 41246 12850
rect 41298 12798 41310 12850
rect 37662 12786 37714 12798
rect 3390 12738 3442 12750
rect 3390 12674 3442 12686
rect 6302 12738 6354 12750
rect 6302 12674 6354 12686
rect 6750 12738 6802 12750
rect 6750 12674 6802 12686
rect 7198 12738 7250 12750
rect 7198 12674 7250 12686
rect 13582 12738 13634 12750
rect 13582 12674 13634 12686
rect 15262 12738 15314 12750
rect 15262 12674 15314 12686
rect 16158 12738 16210 12750
rect 16158 12674 16210 12686
rect 26462 12738 26514 12750
rect 26462 12674 26514 12686
rect 29262 12738 29314 12750
rect 29262 12674 29314 12686
rect 30830 12738 30882 12750
rect 35534 12738 35586 12750
rect 45838 12738 45890 12750
rect 34962 12686 34974 12738
rect 35026 12686 35038 12738
rect 41346 12686 41358 12738
rect 41410 12686 41422 12738
rect 30830 12674 30882 12686
rect 35534 12674 35586 12686
rect 45838 12674 45890 12686
rect 46062 12738 46114 12750
rect 46062 12674 46114 12686
rect 47518 12738 47570 12750
rect 47518 12674 47570 12686
rect 48638 12738 48690 12750
rect 48638 12674 48690 12686
rect 49870 12738 49922 12750
rect 50769 12738 50815 13137
rect 53118 13122 53170 13134
rect 55806 13186 55858 13198
rect 55806 13122 55858 13134
rect 58046 13186 58098 13198
rect 58046 13122 58098 13134
rect 51438 13074 51490 13086
rect 51438 13010 51490 13022
rect 52894 13074 52946 13086
rect 52894 13010 52946 13022
rect 54910 13074 54962 13086
rect 54910 13010 54962 13022
rect 55470 13074 55522 13086
rect 55470 13010 55522 13022
rect 56590 13074 56642 13086
rect 56590 13010 56642 13022
rect 51102 12962 51154 12974
rect 51102 12898 51154 12910
rect 51326 12962 51378 12974
rect 51326 12898 51378 12910
rect 52670 12962 52722 12974
rect 52670 12898 52722 12910
rect 53678 12962 53730 12974
rect 53678 12898 53730 12910
rect 54462 12962 54514 12974
rect 54462 12898 54514 12910
rect 55246 12962 55298 12974
rect 55246 12898 55298 12910
rect 56030 12962 56082 12974
rect 56030 12898 56082 12910
rect 56478 12962 56530 12974
rect 56478 12898 56530 12910
rect 56702 12962 56754 12974
rect 56702 12898 56754 12910
rect 57262 12962 57314 12974
rect 57262 12898 57314 12910
rect 51550 12850 51602 12862
rect 51550 12786 51602 12798
rect 51998 12850 52050 12862
rect 57934 12850 57986 12862
rect 53330 12798 53342 12850
rect 53394 12798 53406 12850
rect 51998 12786 52050 12798
rect 57934 12786 57986 12798
rect 54014 12738 54066 12750
rect 50754 12686 50766 12738
rect 50818 12686 50830 12738
rect 53218 12686 53230 12738
rect 53282 12686 53294 12738
rect 49870 12674 49922 12686
rect 54014 12674 54066 12686
rect 57038 12738 57090 12750
rect 57038 12674 57090 12686
rect 57150 12738 57202 12750
rect 57150 12674 57202 12686
rect 57486 12738 57538 12750
rect 57486 12674 57538 12686
rect 58046 12738 58098 12750
rect 58046 12674 58098 12686
rect 1344 12570 58731 12604
rect 1344 12518 15520 12570
rect 15572 12518 15624 12570
rect 15676 12518 15728 12570
rect 15780 12518 29827 12570
rect 29879 12518 29931 12570
rect 29983 12518 30035 12570
rect 30087 12518 44134 12570
rect 44186 12518 44238 12570
rect 44290 12518 44342 12570
rect 44394 12518 58441 12570
rect 58493 12518 58545 12570
rect 58597 12518 58649 12570
rect 58701 12518 58731 12570
rect 1344 12484 58731 12518
rect 1934 12402 1986 12414
rect 1934 12338 1986 12350
rect 9662 12402 9714 12414
rect 9662 12338 9714 12350
rect 10558 12402 10610 12414
rect 10558 12338 10610 12350
rect 11006 12402 11058 12414
rect 11006 12338 11058 12350
rect 11454 12402 11506 12414
rect 14142 12402 14194 12414
rect 12786 12350 12798 12402
rect 12850 12350 12862 12402
rect 11454 12338 11506 12350
rect 14142 12338 14194 12350
rect 15822 12402 15874 12414
rect 15822 12338 15874 12350
rect 16382 12402 16434 12414
rect 16382 12338 16434 12350
rect 18510 12402 18562 12414
rect 18510 12338 18562 12350
rect 18734 12402 18786 12414
rect 18734 12338 18786 12350
rect 18846 12402 18898 12414
rect 18846 12338 18898 12350
rect 19630 12402 19682 12414
rect 19630 12338 19682 12350
rect 22094 12402 22146 12414
rect 22094 12338 22146 12350
rect 22542 12402 22594 12414
rect 22542 12338 22594 12350
rect 22990 12402 23042 12414
rect 22990 12338 23042 12350
rect 24670 12402 24722 12414
rect 24670 12338 24722 12350
rect 29150 12402 29202 12414
rect 29150 12338 29202 12350
rect 31278 12402 31330 12414
rect 31278 12338 31330 12350
rect 36766 12402 36818 12414
rect 36766 12338 36818 12350
rect 44382 12402 44434 12414
rect 44382 12338 44434 12350
rect 45614 12402 45666 12414
rect 45614 12338 45666 12350
rect 47518 12402 47570 12414
rect 47518 12338 47570 12350
rect 47854 12402 47906 12414
rect 47854 12338 47906 12350
rect 48078 12402 48130 12414
rect 48078 12338 48130 12350
rect 50094 12402 50146 12414
rect 50094 12338 50146 12350
rect 50766 12402 50818 12414
rect 50766 12338 50818 12350
rect 52558 12402 52610 12414
rect 52558 12338 52610 12350
rect 53006 12402 53058 12414
rect 53006 12338 53058 12350
rect 55358 12402 55410 12414
rect 55358 12338 55410 12350
rect 55582 12402 55634 12414
rect 55582 12338 55634 12350
rect 55806 12402 55858 12414
rect 55806 12338 55858 12350
rect 57598 12402 57650 12414
rect 57598 12338 57650 12350
rect 5630 12290 5682 12302
rect 18398 12290 18450 12302
rect 2818 12238 2830 12290
rect 2882 12238 2894 12290
rect 3826 12238 3838 12290
rect 3890 12238 3902 12290
rect 6178 12238 6190 12290
rect 6242 12238 6254 12290
rect 15026 12238 15038 12290
rect 15090 12238 15102 12290
rect 5630 12226 5682 12238
rect 18398 12226 18450 12238
rect 19070 12290 19122 12302
rect 19070 12226 19122 12238
rect 31054 12290 31106 12302
rect 47742 12290 47794 12302
rect 35074 12238 35086 12290
rect 35138 12238 35150 12290
rect 37426 12238 37438 12290
rect 37490 12238 37502 12290
rect 31054 12226 31106 12238
rect 47742 12226 47794 12238
rect 49646 12290 49698 12302
rect 49646 12226 49698 12238
rect 51326 12290 51378 12302
rect 51326 12226 51378 12238
rect 51662 12290 51714 12302
rect 51662 12226 51714 12238
rect 52110 12290 52162 12302
rect 52110 12226 52162 12238
rect 55694 12290 55746 12302
rect 55694 12226 55746 12238
rect 57710 12290 57762 12302
rect 57710 12226 57762 12238
rect 19182 12178 19234 12190
rect 1586 12126 1598 12178
rect 1650 12175 1662 12178
rect 1810 12175 1822 12178
rect 1650 12129 1822 12175
rect 1650 12126 1662 12129
rect 1810 12126 1822 12129
rect 1874 12126 1886 12178
rect 2482 12126 2494 12178
rect 2546 12126 2558 12178
rect 3938 12126 3950 12178
rect 4002 12126 4014 12178
rect 6962 12126 6974 12178
rect 7026 12126 7038 12178
rect 12226 12126 12238 12178
rect 12290 12126 12302 12178
rect 12562 12126 12574 12178
rect 12626 12126 12638 12178
rect 14914 12126 14926 12178
rect 14978 12126 14990 12178
rect 19182 12114 19234 12126
rect 23326 12178 23378 12190
rect 29486 12178 29538 12190
rect 45166 12178 45218 12190
rect 23538 12126 23550 12178
rect 23602 12126 23614 12178
rect 25554 12126 25566 12178
rect 25618 12126 25630 12178
rect 26114 12126 26126 12178
rect 26178 12126 26190 12178
rect 28130 12126 28142 12178
rect 28194 12126 28206 12178
rect 28354 12126 28366 12178
rect 28418 12126 28430 12178
rect 34178 12126 34190 12178
rect 34242 12126 34254 12178
rect 35858 12126 35870 12178
rect 35922 12126 35934 12178
rect 37986 12126 37998 12178
rect 38050 12126 38062 12178
rect 41794 12126 41806 12178
rect 41858 12126 41870 12178
rect 23326 12114 23378 12126
rect 29486 12114 29538 12126
rect 45166 12114 45218 12126
rect 48862 12178 48914 12190
rect 48862 12114 48914 12126
rect 49422 12178 49474 12190
rect 49422 12114 49474 12126
rect 51102 12178 51154 12190
rect 51102 12114 51154 12126
rect 54238 12178 54290 12190
rect 54238 12114 54290 12126
rect 54686 12178 54738 12190
rect 54686 12114 54738 12126
rect 54798 12178 54850 12190
rect 54798 12114 54850 12126
rect 54910 12178 54962 12190
rect 54910 12114 54962 12126
rect 56702 12178 56754 12190
rect 56702 12114 56754 12126
rect 57150 12178 57202 12190
rect 57150 12114 57202 12126
rect 57374 12178 57426 12190
rect 57922 12126 57934 12178
rect 57986 12126 57998 12178
rect 58146 12126 58158 12178
rect 58210 12126 58222 12178
rect 57374 12114 57426 12126
rect 8094 12066 8146 12078
rect 8094 12002 8146 12014
rect 8542 12066 8594 12078
rect 8542 12002 8594 12014
rect 8990 12066 9042 12078
rect 8990 12002 9042 12014
rect 10110 12066 10162 12078
rect 13694 12066 13746 12078
rect 12002 12014 12014 12066
rect 12066 12014 12078 12066
rect 10110 12002 10162 12014
rect 13694 12002 13746 12014
rect 17614 12066 17666 12078
rect 17614 12002 17666 12014
rect 18062 12066 18114 12078
rect 18062 12002 18114 12014
rect 21646 12066 21698 12078
rect 21646 12002 21698 12014
rect 24110 12066 24162 12078
rect 31166 12066 31218 12078
rect 44718 12066 44770 12078
rect 27346 12014 27358 12066
rect 27410 12014 27422 12066
rect 27906 12014 27918 12066
rect 27970 12014 27982 12066
rect 42018 12014 42030 12066
rect 42082 12014 42094 12066
rect 43026 12014 43038 12066
rect 43090 12014 43102 12066
rect 24110 12002 24162 12014
rect 31166 12002 31218 12014
rect 44718 12002 44770 12014
rect 46958 12066 47010 12078
rect 51550 12066 51602 12078
rect 49298 12014 49310 12066
rect 49362 12014 49374 12066
rect 46958 12002 47010 12014
rect 51550 12002 51602 12014
rect 53790 12066 53842 12078
rect 53790 12002 53842 12014
rect 57262 12066 57314 12078
rect 57262 12002 57314 12014
rect 14478 11954 14530 11966
rect 7298 11902 7310 11954
rect 7362 11902 7374 11954
rect 14478 11890 14530 11902
rect 44942 11954 44994 11966
rect 44942 11890 44994 11902
rect 49086 11954 49138 11966
rect 49086 11890 49138 11902
rect 1344 11786 58576 11820
rect 1344 11734 8367 11786
rect 8419 11734 8471 11786
rect 8523 11734 8575 11786
rect 8627 11734 22674 11786
rect 22726 11734 22778 11786
rect 22830 11734 22882 11786
rect 22934 11734 36981 11786
rect 37033 11734 37085 11786
rect 37137 11734 37189 11786
rect 37241 11734 51288 11786
rect 51340 11734 51392 11786
rect 51444 11734 51496 11786
rect 51548 11734 58576 11786
rect 1344 11700 58576 11734
rect 2270 11618 2322 11630
rect 2270 11554 2322 11566
rect 2718 11618 2770 11630
rect 9662 11618 9714 11630
rect 6962 11566 6974 11618
rect 7026 11566 7038 11618
rect 2718 11554 2770 11566
rect 9662 11554 9714 11566
rect 11790 11618 11842 11630
rect 11790 11554 11842 11566
rect 21870 11618 21922 11630
rect 21870 11554 21922 11566
rect 22094 11618 22146 11630
rect 22094 11554 22146 11566
rect 30158 11618 30210 11630
rect 30158 11554 30210 11566
rect 4510 11506 4562 11518
rect 4510 11442 4562 11454
rect 4958 11506 5010 11518
rect 4958 11442 5010 11454
rect 5742 11506 5794 11518
rect 5742 11442 5794 11454
rect 10782 11506 10834 11518
rect 10782 11442 10834 11454
rect 11230 11506 11282 11518
rect 11230 11442 11282 11454
rect 12574 11506 12626 11518
rect 12574 11442 12626 11454
rect 13022 11506 13074 11518
rect 13022 11442 13074 11454
rect 13694 11506 13746 11518
rect 13694 11442 13746 11454
rect 14142 11506 14194 11518
rect 14142 11442 14194 11454
rect 14590 11506 14642 11518
rect 14590 11442 14642 11454
rect 18958 11506 19010 11518
rect 18958 11442 19010 11454
rect 26238 11506 26290 11518
rect 26238 11442 26290 11454
rect 26798 11506 26850 11518
rect 26798 11442 26850 11454
rect 31166 11506 31218 11518
rect 40014 11506 40066 11518
rect 44942 11506 44994 11518
rect 39442 11454 39454 11506
rect 39506 11454 39518 11506
rect 41906 11454 41918 11506
rect 41970 11454 41982 11506
rect 31166 11442 31218 11454
rect 40014 11442 40066 11454
rect 44942 11442 44994 11454
rect 45950 11506 46002 11518
rect 45950 11442 46002 11454
rect 47518 11506 47570 11518
rect 47518 11442 47570 11454
rect 48302 11506 48354 11518
rect 48302 11442 48354 11454
rect 49086 11506 49138 11518
rect 49086 11442 49138 11454
rect 50318 11506 50370 11518
rect 50318 11442 50370 11454
rect 50654 11506 50706 11518
rect 53566 11506 53618 11518
rect 51762 11454 51774 11506
rect 51826 11454 51838 11506
rect 50654 11442 50706 11454
rect 53566 11442 53618 11454
rect 54014 11506 54066 11518
rect 54014 11442 54066 11454
rect 57486 11506 57538 11518
rect 57486 11442 57538 11454
rect 2494 11394 2546 11406
rect 7870 11394 7922 11406
rect 6850 11342 6862 11394
rect 6914 11342 6926 11394
rect 2494 11330 2546 11342
rect 7870 11330 7922 11342
rect 9438 11394 9490 11406
rect 20750 11394 20802 11406
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 19282 11342 19294 11394
rect 19346 11342 19358 11394
rect 9438 11330 9490 11342
rect 20750 11330 20802 11342
rect 22318 11394 22370 11406
rect 22318 11330 22370 11342
rect 23326 11394 23378 11406
rect 30382 11394 30434 11406
rect 44718 11394 44770 11406
rect 23762 11342 23774 11394
rect 23826 11342 23838 11394
rect 23986 11342 23998 11394
rect 24050 11342 24062 11394
rect 27122 11342 27134 11394
rect 27186 11342 27198 11394
rect 38658 11342 38670 11394
rect 38722 11342 38734 11394
rect 38994 11342 39006 11394
rect 39058 11342 39070 11394
rect 40226 11342 40238 11394
rect 40290 11342 40302 11394
rect 41682 11342 41694 11394
rect 41746 11342 41758 11394
rect 23326 11330 23378 11342
rect 30382 11330 30434 11342
rect 44718 11330 44770 11342
rect 45278 11394 45330 11406
rect 55134 11394 55186 11406
rect 51650 11342 51662 11394
rect 51714 11342 51726 11394
rect 45278 11330 45330 11342
rect 55134 11330 55186 11342
rect 55918 11394 55970 11406
rect 55918 11330 55970 11342
rect 56254 11394 56306 11406
rect 56254 11330 56306 11342
rect 56702 11394 56754 11406
rect 56702 11330 56754 11342
rect 2046 11282 2098 11294
rect 15262 11282 15314 11294
rect 7074 11230 7086 11282
rect 7138 11230 7150 11282
rect 9090 11230 9102 11282
rect 9154 11230 9166 11282
rect 2046 11218 2098 11230
rect 15262 11218 15314 11230
rect 19630 11282 19682 11294
rect 19630 11218 19682 11230
rect 22542 11282 22594 11294
rect 22542 11218 22594 11230
rect 22990 11282 23042 11294
rect 22990 11218 23042 11230
rect 23102 11282 23154 11294
rect 30046 11282 30098 11294
rect 33182 11282 33234 11294
rect 25778 11230 25790 11282
rect 25842 11230 25854 11282
rect 28130 11230 28142 11282
rect 28194 11230 28206 11282
rect 31266 11230 31278 11282
rect 31330 11230 31342 11282
rect 32946 11230 32958 11282
rect 33010 11230 33022 11282
rect 23102 11218 23154 11230
rect 30046 11218 30098 11230
rect 33182 11218 33234 11230
rect 39902 11282 39954 11294
rect 39902 11218 39954 11230
rect 44270 11282 44322 11294
rect 44270 11218 44322 11230
rect 45166 11282 45218 11294
rect 45166 11218 45218 11230
rect 46846 11282 46898 11294
rect 46846 11218 46898 11230
rect 46958 11282 47010 11294
rect 46958 11218 47010 11230
rect 52110 11282 52162 11294
rect 52110 11218 52162 11230
rect 54910 11282 54962 11294
rect 54910 11218 54962 11230
rect 57822 11282 57874 11294
rect 57822 11218 57874 11230
rect 3166 11170 3218 11182
rect 3166 11106 3218 11118
rect 3502 11170 3554 11182
rect 3502 11106 3554 11118
rect 3950 11170 4002 11182
rect 3950 11106 4002 11118
rect 6190 11170 6242 11182
rect 11678 11170 11730 11182
rect 9986 11118 9998 11170
rect 10050 11118 10062 11170
rect 6190 11106 6242 11118
rect 11678 11106 11730 11118
rect 15710 11170 15762 11182
rect 15710 11106 15762 11118
rect 19518 11170 19570 11182
rect 19518 11106 19570 11118
rect 21422 11170 21474 11182
rect 29822 11170 29874 11182
rect 28466 11118 28478 11170
rect 28530 11118 28542 11170
rect 21422 11106 21474 11118
rect 29822 11106 29874 11118
rect 38222 11170 38274 11182
rect 38222 11106 38274 11118
rect 40686 11170 40738 11182
rect 40686 11106 40738 11118
rect 42926 11170 42978 11182
rect 42926 11106 42978 11118
rect 46286 11170 46338 11182
rect 46286 11106 46338 11118
rect 47182 11170 47234 11182
rect 47182 11106 47234 11118
rect 48638 11170 48690 11182
rect 48638 11106 48690 11118
rect 49534 11170 49586 11182
rect 49534 11106 49586 11118
rect 54686 11170 54738 11182
rect 56366 11170 56418 11182
rect 55458 11118 55470 11170
rect 55522 11118 55534 11170
rect 54686 11106 54738 11118
rect 56366 11106 56418 11118
rect 57374 11170 57426 11182
rect 57374 11106 57426 11118
rect 57598 11170 57650 11182
rect 57598 11106 57650 11118
rect 1344 11002 58731 11036
rect 1344 10950 15520 11002
rect 15572 10950 15624 11002
rect 15676 10950 15728 11002
rect 15780 10950 29827 11002
rect 29879 10950 29931 11002
rect 29983 10950 30035 11002
rect 30087 10950 44134 11002
rect 44186 10950 44238 11002
rect 44290 10950 44342 11002
rect 44394 10950 58441 11002
rect 58493 10950 58545 11002
rect 58597 10950 58649 11002
rect 58701 10950 58731 11002
rect 1344 10916 58731 10950
rect 2270 10834 2322 10846
rect 2270 10770 2322 10782
rect 15486 10834 15538 10846
rect 15486 10770 15538 10782
rect 24110 10834 24162 10846
rect 24110 10770 24162 10782
rect 24670 10834 24722 10846
rect 24670 10770 24722 10782
rect 25902 10834 25954 10846
rect 25902 10770 25954 10782
rect 26574 10834 26626 10846
rect 26574 10770 26626 10782
rect 27358 10834 27410 10846
rect 27358 10770 27410 10782
rect 29150 10834 29202 10846
rect 29150 10770 29202 10782
rect 29934 10834 29986 10846
rect 29934 10770 29986 10782
rect 30494 10834 30546 10846
rect 30494 10770 30546 10782
rect 38334 10834 38386 10846
rect 38334 10770 38386 10782
rect 55246 10834 55298 10846
rect 55246 10770 55298 10782
rect 55806 10834 55858 10846
rect 55806 10770 55858 10782
rect 56030 10834 56082 10846
rect 56030 10770 56082 10782
rect 56142 10834 56194 10846
rect 56142 10770 56194 10782
rect 9662 10722 9714 10734
rect 13470 10722 13522 10734
rect 3042 10670 3054 10722
rect 3106 10670 3118 10722
rect 12114 10670 12126 10722
rect 12178 10670 12190 10722
rect 12562 10670 12574 10722
rect 12626 10670 12638 10722
rect 9662 10658 9714 10670
rect 13470 10658 13522 10670
rect 13582 10722 13634 10734
rect 13582 10658 13634 10670
rect 14142 10722 14194 10734
rect 14142 10658 14194 10670
rect 16606 10722 16658 10734
rect 16606 10658 16658 10670
rect 17390 10722 17442 10734
rect 21646 10722 21698 10734
rect 19282 10670 19294 10722
rect 19346 10670 19358 10722
rect 17390 10658 17442 10670
rect 21646 10658 21698 10670
rect 21870 10722 21922 10734
rect 21870 10658 21922 10670
rect 29486 10722 29538 10734
rect 29486 10658 29538 10670
rect 32286 10722 32338 10734
rect 39342 10722 39394 10734
rect 34962 10670 34974 10722
rect 35026 10670 35038 10722
rect 36306 10670 36318 10722
rect 36370 10670 36382 10722
rect 32286 10658 32338 10670
rect 39342 10658 39394 10670
rect 40014 10722 40066 10734
rect 42030 10722 42082 10734
rect 41234 10670 41246 10722
rect 41298 10670 41310 10722
rect 40014 10658 40066 10670
rect 42030 10658 42082 10670
rect 46398 10722 46450 10734
rect 46398 10658 46450 10670
rect 46622 10722 46674 10734
rect 46622 10658 46674 10670
rect 47294 10722 47346 10734
rect 47294 10658 47346 10670
rect 48862 10722 48914 10734
rect 48862 10658 48914 10670
rect 49758 10722 49810 10734
rect 49758 10658 49810 10670
rect 49982 10722 50034 10734
rect 55582 10722 55634 10734
rect 51762 10670 51774 10722
rect 51826 10670 51838 10722
rect 49982 10658 50034 10670
rect 55582 10658 55634 10670
rect 10670 10610 10722 10622
rect 13022 10610 13074 10622
rect 2930 10558 2942 10610
rect 2994 10558 3006 10610
rect 5618 10558 5630 10610
rect 5682 10558 5694 10610
rect 7186 10558 7198 10610
rect 7250 10558 7262 10610
rect 7410 10558 7422 10610
rect 7474 10558 7486 10610
rect 11218 10558 11230 10610
rect 11282 10558 11294 10610
rect 10670 10546 10722 10558
rect 13022 10546 13074 10558
rect 14366 10610 14418 10622
rect 14366 10546 14418 10558
rect 14590 10610 14642 10622
rect 14590 10546 14642 10558
rect 14702 10610 14754 10622
rect 14702 10546 14754 10558
rect 15374 10610 15426 10622
rect 15374 10546 15426 10558
rect 15710 10610 15762 10622
rect 15710 10546 15762 10558
rect 16270 10610 16322 10622
rect 16270 10546 16322 10558
rect 17614 10610 17666 10622
rect 21086 10610 21138 10622
rect 23326 10610 23378 10622
rect 20738 10558 20750 10610
rect 20802 10558 20814 10610
rect 22418 10558 22430 10610
rect 22482 10558 22494 10610
rect 22866 10558 22878 10610
rect 22930 10558 22942 10610
rect 17614 10546 17666 10558
rect 21086 10546 21138 10558
rect 23326 10546 23378 10558
rect 25454 10610 25506 10622
rect 25454 10546 25506 10558
rect 26350 10610 26402 10622
rect 26350 10546 26402 10558
rect 26574 10610 26626 10622
rect 26574 10546 26626 10558
rect 26910 10610 26962 10622
rect 31502 10610 31554 10622
rect 39118 10610 39170 10622
rect 28130 10558 28142 10610
rect 28194 10558 28206 10610
rect 28354 10558 28366 10610
rect 28418 10558 28430 10610
rect 31714 10558 31726 10610
rect 31778 10558 31790 10610
rect 34850 10558 34862 10610
rect 34914 10558 34926 10610
rect 26910 10546 26962 10558
rect 31502 10546 31554 10558
rect 39118 10546 39170 10558
rect 39566 10610 39618 10622
rect 39566 10546 39618 10558
rect 40126 10610 40178 10622
rect 41918 10610 41970 10622
rect 41570 10558 41582 10610
rect 41634 10558 41646 10610
rect 40126 10546 40178 10558
rect 41918 10546 41970 10558
rect 42254 10610 42306 10622
rect 42254 10546 42306 10558
rect 43038 10610 43090 10622
rect 47406 10610 47458 10622
rect 43474 10558 43486 10610
rect 43538 10558 43550 10610
rect 45042 10558 45054 10610
rect 45106 10558 45118 10610
rect 43038 10546 43090 10558
rect 47406 10546 47458 10558
rect 47854 10610 47906 10622
rect 47854 10546 47906 10558
rect 49310 10610 49362 10622
rect 51986 10558 51998 10610
rect 52050 10558 52062 10610
rect 52882 10558 52894 10610
rect 52946 10558 52958 10610
rect 56914 10558 56926 10610
rect 56978 10558 56990 10610
rect 49310 10546 49362 10558
rect 13806 10498 13858 10510
rect 3042 10446 3054 10498
rect 3106 10446 3118 10498
rect 4946 10446 4958 10498
rect 5010 10446 5022 10498
rect 5842 10446 5854 10498
rect 5906 10446 5918 10498
rect 13806 10434 13858 10446
rect 14478 10498 14530 10510
rect 39790 10498 39842 10510
rect 49534 10498 49586 10510
rect 28802 10446 28814 10498
rect 28866 10446 28878 10498
rect 40898 10446 40910 10498
rect 40962 10446 40974 10498
rect 45266 10446 45278 10498
rect 45330 10446 45342 10498
rect 46722 10446 46734 10498
rect 46786 10446 46798 10498
rect 47618 10446 47630 10498
rect 47682 10446 47694 10498
rect 14478 10434 14530 10446
rect 39790 10434 39842 10446
rect 49534 10434 49586 10446
rect 50430 10498 50482 10510
rect 50430 10434 50482 10446
rect 54686 10498 54738 10510
rect 54686 10434 54738 10446
rect 9886 10386 9938 10398
rect 10782 10386 10834 10398
rect 2818 10334 2830 10386
rect 2882 10334 2894 10386
rect 8306 10334 8318 10386
rect 8370 10334 8382 10386
rect 10210 10334 10222 10386
rect 10274 10334 10286 10386
rect 9886 10322 9938 10334
rect 10782 10322 10834 10334
rect 12798 10386 12850 10398
rect 12798 10322 12850 10334
rect 16046 10386 16098 10398
rect 16046 10322 16098 10334
rect 16718 10386 16770 10398
rect 16718 10322 16770 10334
rect 16830 10386 16882 10398
rect 16830 10322 16882 10334
rect 17838 10386 17890 10398
rect 17838 10322 17890 10334
rect 18062 10386 18114 10398
rect 18062 10322 18114 10334
rect 18510 10386 18562 10398
rect 18510 10322 18562 10334
rect 21982 10386 22034 10398
rect 29374 10386 29426 10398
rect 23426 10334 23438 10386
rect 23490 10334 23502 10386
rect 21982 10322 22034 10334
rect 29374 10322 29426 10334
rect 37662 10386 37714 10398
rect 48078 10386 48130 10398
rect 38770 10334 38782 10386
rect 38834 10334 38846 10386
rect 37662 10322 37714 10334
rect 48078 10322 48130 10334
rect 54238 10386 54290 10398
rect 57934 10386 57986 10398
rect 54674 10334 54686 10386
rect 54738 10383 54750 10386
rect 55122 10383 55134 10386
rect 54738 10337 55134 10383
rect 54738 10334 54750 10337
rect 55122 10334 55134 10337
rect 55186 10334 55198 10386
rect 54238 10322 54290 10334
rect 57934 10322 57986 10334
rect 1344 10218 58576 10252
rect 1344 10166 8367 10218
rect 8419 10166 8471 10218
rect 8523 10166 8575 10218
rect 8627 10166 22674 10218
rect 22726 10166 22778 10218
rect 22830 10166 22882 10218
rect 22934 10166 36981 10218
rect 37033 10166 37085 10218
rect 37137 10166 37189 10218
rect 37241 10166 51288 10218
rect 51340 10166 51392 10218
rect 51444 10166 51496 10218
rect 51548 10166 58576 10218
rect 1344 10132 58576 10166
rect 13918 10050 13970 10062
rect 47966 10050 48018 10062
rect 4610 9998 4622 10050
rect 4674 9998 4686 10050
rect 6626 9998 6638 10050
rect 6690 9998 6702 10050
rect 9426 9998 9438 10050
rect 9490 9998 9502 10050
rect 19954 9998 19966 10050
rect 20018 9998 20030 10050
rect 27010 9998 27022 10050
rect 27074 10047 27086 10050
rect 28018 10047 28030 10050
rect 27074 10001 28030 10047
rect 27074 9998 27086 10001
rect 28018 9998 28030 10001
rect 28082 9998 28094 10050
rect 13918 9986 13970 9998
rect 47966 9986 48018 9998
rect 49646 10050 49698 10062
rect 49646 9986 49698 9998
rect 11566 9938 11618 9950
rect 4498 9886 4510 9938
rect 4562 9886 4574 9938
rect 6738 9886 6750 9938
rect 6802 9886 6814 9938
rect 11566 9874 11618 9886
rect 13694 9938 13746 9950
rect 13694 9874 13746 9886
rect 14254 9938 14306 9950
rect 18286 9938 18338 9950
rect 15362 9886 15374 9938
rect 15426 9886 15438 9938
rect 14254 9874 14306 9886
rect 18286 9874 18338 9886
rect 27582 9938 27634 9950
rect 27582 9874 27634 9886
rect 28030 9938 28082 9950
rect 28030 9874 28082 9886
rect 30718 9938 30770 9950
rect 30718 9874 30770 9886
rect 38446 9938 38498 9950
rect 49982 9938 50034 9950
rect 41794 9886 41806 9938
rect 41858 9886 41870 9938
rect 42914 9886 42926 9938
rect 42978 9886 42990 9938
rect 46946 9886 46958 9938
rect 47010 9886 47022 9938
rect 38446 9874 38498 9886
rect 49982 9874 50034 9886
rect 3950 9826 4002 9838
rect 9102 9826 9154 9838
rect 1922 9774 1934 9826
rect 1986 9774 1998 9826
rect 4162 9774 4174 9826
rect 4226 9774 4238 9826
rect 6066 9774 6078 9826
rect 6130 9774 6142 9826
rect 6290 9774 6302 9826
rect 6354 9774 6366 9826
rect 7634 9774 7646 9826
rect 7698 9774 7710 9826
rect 3950 9762 4002 9774
rect 9102 9762 9154 9774
rect 9998 9826 10050 9838
rect 9998 9762 10050 9774
rect 10446 9826 10498 9838
rect 16158 9826 16210 9838
rect 42590 9826 42642 9838
rect 15698 9774 15710 9826
rect 15762 9774 15774 9826
rect 18946 9774 18958 9826
rect 19010 9774 19022 9826
rect 22642 9774 22654 9826
rect 22706 9774 22718 9826
rect 24658 9774 24670 9826
rect 24722 9774 24734 9826
rect 30258 9774 30270 9826
rect 30322 9774 30334 9826
rect 31266 9774 31278 9826
rect 31330 9774 31342 9826
rect 31602 9774 31614 9826
rect 31666 9774 31678 9826
rect 34290 9774 34302 9826
rect 34354 9774 34366 9826
rect 35186 9774 35198 9826
rect 35250 9774 35262 9826
rect 38098 9774 38110 9826
rect 38162 9774 38174 9826
rect 40114 9774 40126 9826
rect 40178 9774 40190 9826
rect 40450 9774 40462 9826
rect 40514 9774 40526 9826
rect 10446 9762 10498 9774
rect 16158 9762 16210 9774
rect 42590 9762 42642 9774
rect 45054 9826 45106 9838
rect 48190 9826 48242 9838
rect 46722 9774 46734 9826
rect 46786 9774 46798 9826
rect 45054 9762 45106 9774
rect 48190 9762 48242 9774
rect 48414 9826 48466 9838
rect 48414 9762 48466 9774
rect 48526 9826 48578 9838
rect 56030 9826 56082 9838
rect 49074 9774 49086 9826
rect 49138 9774 49150 9826
rect 49298 9774 49310 9826
rect 49362 9774 49374 9826
rect 48526 9762 48578 9774
rect 56030 9762 56082 9774
rect 56478 9826 56530 9838
rect 56478 9762 56530 9774
rect 8878 9714 8930 9726
rect 2482 9662 2494 9714
rect 2546 9662 2558 9714
rect 7746 9662 7758 9714
rect 7810 9662 7822 9714
rect 8878 9650 8930 9662
rect 11230 9714 11282 9726
rect 11230 9650 11282 9662
rect 17838 9714 17890 9726
rect 23214 9714 23266 9726
rect 38334 9714 38386 9726
rect 42366 9714 42418 9726
rect 49534 9714 49586 9726
rect 18834 9662 18846 9714
rect 18898 9662 18910 9714
rect 26338 9662 26350 9714
rect 26402 9662 26414 9714
rect 32834 9662 32846 9714
rect 32898 9662 32910 9714
rect 34178 9662 34190 9714
rect 34242 9662 34254 9714
rect 36418 9662 36430 9714
rect 36482 9662 36494 9714
rect 39330 9662 39342 9714
rect 39394 9662 39406 9714
rect 40338 9662 40350 9714
rect 40402 9662 40414 9714
rect 46498 9662 46510 9714
rect 46562 9662 46574 9714
rect 17838 9650 17890 9662
rect 23214 9650 23266 9662
rect 38334 9650 38386 9662
rect 42366 9650 42418 9662
rect 49534 9650 49586 9662
rect 54910 9714 54962 9726
rect 58146 9662 58158 9714
rect 58210 9662 58222 9714
rect 54910 9650 54962 9662
rect 12574 9602 12626 9614
rect 8082 9550 8094 9602
rect 8146 9550 8158 9602
rect 12574 9538 12626 9550
rect 14702 9602 14754 9614
rect 27022 9602 27074 9614
rect 24098 9550 24110 9602
rect 24162 9550 24174 9602
rect 14702 9538 14754 9550
rect 27022 9538 27074 9550
rect 30606 9602 30658 9614
rect 30606 9538 30658 9550
rect 30830 9602 30882 9614
rect 30830 9538 30882 9550
rect 42814 9602 42866 9614
rect 42814 9538 42866 9550
rect 42926 9602 42978 9614
rect 42926 9538 42978 9550
rect 43486 9602 43538 9614
rect 43486 9538 43538 9550
rect 48078 9602 48130 9614
rect 54562 9550 54574 9602
rect 54626 9550 54638 9602
rect 48078 9538 48130 9550
rect 1344 9434 58731 9468
rect 1344 9382 15520 9434
rect 15572 9382 15624 9434
rect 15676 9382 15728 9434
rect 15780 9382 29827 9434
rect 29879 9382 29931 9434
rect 29983 9382 30035 9434
rect 30087 9382 44134 9434
rect 44186 9382 44238 9434
rect 44290 9382 44342 9434
rect 44394 9382 58441 9434
rect 58493 9382 58545 9434
rect 58597 9382 58649 9434
rect 58701 9382 58731 9434
rect 1344 9348 58731 9382
rect 5070 9266 5122 9278
rect 5070 9202 5122 9214
rect 7534 9266 7586 9278
rect 7534 9202 7586 9214
rect 7982 9266 8034 9278
rect 7982 9202 8034 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 10110 9266 10162 9278
rect 10110 9202 10162 9214
rect 21646 9266 21698 9278
rect 21646 9202 21698 9214
rect 39454 9266 39506 9278
rect 47070 9266 47122 9278
rect 41010 9214 41022 9266
rect 41074 9214 41086 9266
rect 39454 9202 39506 9214
rect 47070 9202 47122 9214
rect 50430 9266 50482 9278
rect 50430 9202 50482 9214
rect 3726 9154 3778 9166
rect 3726 9090 3778 9102
rect 3838 9154 3890 9166
rect 3838 9090 3890 9102
rect 4510 9154 4562 9166
rect 4510 9090 4562 9102
rect 4846 9154 4898 9166
rect 4846 9090 4898 9102
rect 5182 9154 5234 9166
rect 5182 9090 5234 9102
rect 7086 9154 7138 9166
rect 7086 9090 7138 9102
rect 10670 9154 10722 9166
rect 10670 9090 10722 9102
rect 11230 9154 11282 9166
rect 11230 9090 11282 9102
rect 13806 9154 13858 9166
rect 15598 9154 15650 9166
rect 14690 9102 14702 9154
rect 14754 9102 14766 9154
rect 13806 9090 13858 9102
rect 15598 9090 15650 9102
rect 17726 9154 17778 9166
rect 17726 9090 17778 9102
rect 18062 9154 18114 9166
rect 18062 9090 18114 9102
rect 19182 9154 19234 9166
rect 26686 9154 26738 9166
rect 37102 9154 37154 9166
rect 22530 9102 22542 9154
rect 22594 9102 22606 9154
rect 24434 9102 24446 9154
rect 24498 9102 24510 9154
rect 25778 9102 25790 9154
rect 25842 9102 25854 9154
rect 27346 9102 27358 9154
rect 27410 9102 27422 9154
rect 19182 9090 19234 9102
rect 26686 9090 26738 9102
rect 37102 9090 37154 9102
rect 37214 9154 37266 9166
rect 42590 9154 42642 9166
rect 46398 9154 46450 9166
rect 41570 9102 41582 9154
rect 41634 9102 41646 9154
rect 43586 9102 43598 9154
rect 43650 9102 43662 9154
rect 44594 9102 44606 9154
rect 44658 9102 44670 9154
rect 37214 9090 37266 9102
rect 42590 9090 42642 9102
rect 46398 9090 46450 9102
rect 48750 9154 48802 9166
rect 48750 9090 48802 9102
rect 48974 9154 49026 9166
rect 57362 9102 57374 9154
rect 57426 9102 57438 9154
rect 48974 9090 49026 9102
rect 4062 9042 4114 9054
rect 2706 8990 2718 9042
rect 2770 8990 2782 9042
rect 3378 8990 3390 9042
rect 3442 8990 3454 9042
rect 4062 8978 4114 8990
rect 4398 9042 4450 9054
rect 4398 8978 4450 8990
rect 9998 9042 10050 9054
rect 9998 8978 10050 8990
rect 10334 9042 10386 9054
rect 10334 8978 10386 8990
rect 10782 9042 10834 9054
rect 18286 9042 18338 9054
rect 14466 8990 14478 9042
rect 14530 8990 14542 9042
rect 10782 8978 10834 8990
rect 18286 8978 18338 8990
rect 18510 9042 18562 9054
rect 19070 9042 19122 9054
rect 25230 9042 25282 9054
rect 18722 8990 18734 9042
rect 18786 8990 18798 9042
rect 21970 8990 21982 9042
rect 22034 8990 22046 9042
rect 23650 8990 23662 9042
rect 23714 8990 23726 9042
rect 18510 8978 18562 8990
rect 19070 8978 19122 8990
rect 25230 8978 25282 8990
rect 25454 9042 25506 9054
rect 25454 8978 25506 8990
rect 26014 9042 26066 9054
rect 26014 8978 26066 8990
rect 26462 9042 26514 9054
rect 28030 9042 28082 9054
rect 47630 9042 47682 9054
rect 27570 8990 27582 9042
rect 27634 8990 27646 9042
rect 41122 8990 41134 9042
rect 41186 8990 41198 9042
rect 41906 8990 41918 9042
rect 41970 8990 41982 9042
rect 43026 8990 43038 9042
rect 43090 8990 43102 9042
rect 44706 8990 44718 9042
rect 44770 8990 44782 9042
rect 26462 8978 26514 8990
rect 28030 8978 28082 8990
rect 47630 8978 47682 8990
rect 48078 9042 48130 9054
rect 48078 8978 48130 8990
rect 48190 9042 48242 9054
rect 48190 8978 48242 8990
rect 50766 9042 50818 9054
rect 50766 8978 50818 8990
rect 50990 9042 51042 9054
rect 50990 8978 51042 8990
rect 52894 9042 52946 9054
rect 52894 8978 52946 8990
rect 53230 9042 53282 9054
rect 55346 8990 55358 9042
rect 55410 8990 55422 9042
rect 56466 8990 56478 9042
rect 56530 8990 56542 9042
rect 57586 8990 57598 9042
rect 57650 8990 57662 9042
rect 53230 8978 53282 8990
rect 3950 8930 4002 8942
rect 2034 8878 2046 8930
rect 2098 8878 2110 8930
rect 3950 8866 4002 8878
rect 5742 8930 5794 8942
rect 5742 8866 5794 8878
rect 8542 8930 8594 8942
rect 8542 8866 8594 8878
rect 8990 8930 9042 8942
rect 8990 8866 9042 8878
rect 13358 8930 13410 8942
rect 26574 8930 26626 8942
rect 15138 8878 15150 8930
rect 15202 8878 15214 8930
rect 18610 8878 18622 8930
rect 18674 8878 18686 8930
rect 13358 8866 13410 8878
rect 26574 8866 26626 8878
rect 31054 8930 31106 8942
rect 52110 8930 52162 8942
rect 57710 8930 57762 8942
rect 51314 8878 51326 8930
rect 51378 8878 51390 8930
rect 53554 8878 53566 8930
rect 53618 8878 53630 8930
rect 55234 8878 55246 8930
rect 55298 8878 55310 8930
rect 31054 8866 31106 8878
rect 52110 8866 52162 8878
rect 57710 8866 57762 8878
rect 4510 8818 4562 8830
rect 6862 8818 6914 8830
rect 10670 8818 10722 8830
rect 6514 8766 6526 8818
rect 6578 8766 6590 8818
rect 7634 8766 7646 8818
rect 7698 8815 7710 8818
rect 8978 8815 8990 8818
rect 7698 8769 8990 8815
rect 7698 8766 7710 8769
rect 8978 8766 8990 8769
rect 9042 8766 9054 8818
rect 4510 8754 4562 8766
rect 6862 8754 6914 8766
rect 10670 8754 10722 8766
rect 28366 8818 28418 8830
rect 28366 8754 28418 8766
rect 37214 8818 37266 8830
rect 37214 8754 37266 8766
rect 47518 8818 47570 8830
rect 47518 8754 47570 8766
rect 47854 8818 47906 8830
rect 47854 8754 47906 8766
rect 49086 8818 49138 8830
rect 49086 8754 49138 8766
rect 1344 8650 58576 8684
rect 1344 8598 8367 8650
rect 8419 8598 8471 8650
rect 8523 8598 8575 8650
rect 8627 8598 22674 8650
rect 22726 8598 22778 8650
rect 22830 8598 22882 8650
rect 22934 8598 36981 8650
rect 37033 8598 37085 8650
rect 37137 8598 37189 8650
rect 37241 8598 51288 8650
rect 51340 8598 51392 8650
rect 51444 8598 51496 8650
rect 51548 8598 58576 8650
rect 1344 8564 58576 8598
rect 25902 8482 25954 8494
rect 10770 8430 10782 8482
rect 10834 8430 10846 8482
rect 25902 8418 25954 8430
rect 35086 8482 35138 8494
rect 35086 8418 35138 8430
rect 37214 8482 37266 8494
rect 43150 8482 43202 8494
rect 39218 8430 39230 8482
rect 39282 8430 39294 8482
rect 37214 8418 37266 8430
rect 43150 8418 43202 8430
rect 47854 8482 47906 8494
rect 47854 8418 47906 8430
rect 48302 8482 48354 8494
rect 48302 8418 48354 8430
rect 2046 8370 2098 8382
rect 2046 8306 2098 8318
rect 3950 8370 4002 8382
rect 3950 8306 4002 8318
rect 4846 8370 4898 8382
rect 4846 8306 4898 8318
rect 5742 8370 5794 8382
rect 12910 8370 12962 8382
rect 10322 8318 10334 8370
rect 10386 8318 10398 8370
rect 11218 8318 11230 8370
rect 11282 8318 11294 8370
rect 5742 8306 5794 8318
rect 12910 8306 12962 8318
rect 14926 8370 14978 8382
rect 21310 8370 21362 8382
rect 31838 8370 31890 8382
rect 20178 8318 20190 8370
rect 20242 8318 20254 8370
rect 24546 8318 24558 8370
rect 24610 8318 24622 8370
rect 14926 8306 14978 8318
rect 21310 8306 21362 8318
rect 31838 8306 31890 8318
rect 33518 8370 33570 8382
rect 37774 8370 37826 8382
rect 37426 8318 37438 8370
rect 37490 8318 37502 8370
rect 33518 8306 33570 8318
rect 37774 8306 37826 8318
rect 42142 8370 42194 8382
rect 42142 8306 42194 8318
rect 45950 8370 46002 8382
rect 45950 8306 46002 8318
rect 49086 8370 49138 8382
rect 49086 8306 49138 8318
rect 50318 8370 50370 8382
rect 57150 8370 57202 8382
rect 50642 8318 50654 8370
rect 50706 8318 50718 8370
rect 56466 8318 56478 8370
rect 56530 8318 56542 8370
rect 50318 8306 50370 8318
rect 57150 8306 57202 8318
rect 6414 8258 6466 8270
rect 9438 8258 9490 8270
rect 3154 8206 3166 8258
rect 3218 8206 3230 8258
rect 7410 8206 7422 8258
rect 7474 8206 7486 8258
rect 7970 8206 7982 8258
rect 8034 8206 8046 8258
rect 8194 8206 8206 8258
rect 8258 8206 8270 8258
rect 6414 8194 6466 8206
rect 9438 8194 9490 8206
rect 9774 8258 9826 8270
rect 12462 8258 12514 8270
rect 13918 8258 13970 8270
rect 21534 8258 21586 8270
rect 26014 8258 26066 8270
rect 10434 8206 10446 8258
rect 10498 8206 10510 8258
rect 11330 8206 11342 8258
rect 11394 8206 11406 8258
rect 13458 8206 13470 8258
rect 13522 8206 13534 8258
rect 19842 8206 19854 8258
rect 19906 8206 19918 8258
rect 21858 8206 21870 8258
rect 21922 8206 21934 8258
rect 22306 8206 22318 8258
rect 22370 8206 22382 8258
rect 22866 8206 22878 8258
rect 22930 8206 22942 8258
rect 24994 8206 25006 8258
rect 25058 8206 25070 8258
rect 9774 8194 9826 8206
rect 12462 8194 12514 8206
rect 13918 8194 13970 8206
rect 21534 8194 21586 8206
rect 26014 8194 26066 8206
rect 26462 8258 26514 8270
rect 26462 8194 26514 8206
rect 26910 8258 26962 8270
rect 26910 8194 26962 8206
rect 27134 8258 27186 8270
rect 28030 8258 28082 8270
rect 27794 8206 27806 8258
rect 27858 8206 27870 8258
rect 27134 8194 27186 8206
rect 28030 8194 28082 8206
rect 29710 8258 29762 8270
rect 29710 8194 29762 8206
rect 31054 8258 31106 8270
rect 31054 8194 31106 8206
rect 32734 8258 32786 8270
rect 32734 8194 32786 8206
rect 33406 8258 33458 8270
rect 33406 8194 33458 8206
rect 34078 8258 34130 8270
rect 34078 8194 34130 8206
rect 35870 8258 35922 8270
rect 35870 8194 35922 8206
rect 37998 8258 38050 8270
rect 42478 8258 42530 8270
rect 48078 8258 48130 8270
rect 39330 8206 39342 8258
rect 39394 8206 39406 8258
rect 40674 8206 40686 8258
rect 40738 8206 40750 8258
rect 41794 8206 41806 8258
rect 41858 8206 41870 8258
rect 42690 8206 42702 8258
rect 42754 8206 42766 8258
rect 43474 8206 43486 8258
rect 43538 8206 43550 8258
rect 45042 8206 45054 8258
rect 45106 8206 45118 8258
rect 46386 8206 46398 8258
rect 46450 8206 46462 8258
rect 47618 8206 47630 8258
rect 47682 8206 47694 8258
rect 37998 8194 38050 8206
rect 42478 8194 42530 8206
rect 48078 8194 48130 8206
rect 48414 8258 48466 8270
rect 48738 8206 48750 8258
rect 48802 8206 48814 8258
rect 50866 8206 50878 8258
rect 50930 8206 50942 8258
rect 53778 8206 53790 8258
rect 53842 8206 53854 8258
rect 54786 8206 54798 8258
rect 54850 8206 54862 8258
rect 57250 8206 57262 8258
rect 57314 8206 57326 8258
rect 57698 8206 57710 8258
rect 57762 8206 57774 8258
rect 48414 8194 48466 8206
rect 2382 8146 2434 8158
rect 2382 8082 2434 8094
rect 6302 8146 6354 8158
rect 14142 8146 14194 8158
rect 6738 8094 6750 8146
rect 6802 8094 6814 8146
rect 7298 8094 7310 8146
rect 7362 8094 7374 8146
rect 8866 8094 8878 8146
rect 8930 8094 8942 8146
rect 9202 8094 9214 8146
rect 9266 8094 9278 8146
rect 6302 8082 6354 8094
rect 14142 8082 14194 8094
rect 15486 8146 15538 8158
rect 15486 8082 15538 8094
rect 15598 8146 15650 8158
rect 20526 8146 20578 8158
rect 25454 8146 25506 8158
rect 15698 8094 15710 8146
rect 15762 8094 15774 8146
rect 23874 8094 23886 8146
rect 23938 8094 23950 8146
rect 15598 8082 15650 8094
rect 20526 8082 20578 8094
rect 25454 8082 25506 8094
rect 27358 8146 27410 8158
rect 27358 8082 27410 8094
rect 27470 8146 27522 8158
rect 27470 8082 27522 8094
rect 28142 8146 28194 8158
rect 29150 8146 29202 8158
rect 28578 8094 28590 8146
rect 28642 8094 28654 8146
rect 28142 8082 28194 8094
rect 29150 8082 29202 8094
rect 29374 8146 29426 8158
rect 29374 8082 29426 8094
rect 31166 8146 31218 8158
rect 31166 8082 31218 8094
rect 31614 8146 31666 8158
rect 31614 8082 31666 8094
rect 32510 8146 32562 8158
rect 32510 8082 32562 8094
rect 33630 8146 33682 8158
rect 33630 8082 33682 8094
rect 34974 8146 35026 8158
rect 34974 8082 35026 8094
rect 35534 8146 35586 8158
rect 35534 8082 35586 8094
rect 37438 8146 37490 8158
rect 46846 8146 46898 8158
rect 42242 8094 42254 8146
rect 42306 8094 42318 8146
rect 43362 8094 43374 8146
rect 43426 8094 43438 8146
rect 44034 8094 44046 8146
rect 44098 8094 44110 8146
rect 44818 8094 44830 8146
rect 44882 8094 44894 8146
rect 45154 8094 45166 8146
rect 45218 8094 45230 8146
rect 37438 8082 37490 8094
rect 46846 8082 46898 8094
rect 51550 8146 51602 8158
rect 54002 8094 54014 8146
rect 54066 8094 54078 8146
rect 54674 8094 54686 8146
rect 54738 8094 54750 8146
rect 51550 8082 51602 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 2718 8034 2770 8046
rect 2718 7970 2770 7982
rect 6078 8034 6130 8046
rect 6078 7970 6130 7982
rect 7646 8034 7698 8046
rect 7646 7970 7698 7982
rect 7758 8034 7810 8046
rect 7758 7970 7810 7982
rect 13694 8034 13746 8046
rect 13694 7970 13746 7982
rect 13806 8034 13858 8046
rect 13806 7970 13858 7982
rect 15262 8034 15314 8046
rect 15262 7970 15314 7982
rect 15374 8034 15426 8046
rect 15374 7970 15426 7982
rect 25902 8034 25954 8046
rect 25902 7970 25954 7982
rect 29598 8034 29650 8046
rect 29598 7970 29650 7982
rect 31390 8034 31442 8046
rect 35086 8034 35138 8046
rect 32162 7982 32174 8034
rect 32226 7982 32238 8034
rect 33058 7982 33070 8034
rect 33122 7982 33134 8034
rect 31390 7970 31442 7982
rect 35086 7970 35138 7982
rect 35646 8034 35698 8046
rect 35646 7970 35698 7982
rect 45838 8034 45890 8046
rect 45838 7970 45890 7982
rect 46062 8034 46114 8046
rect 46062 7970 46114 7982
rect 46734 8034 46786 8046
rect 46734 7970 46786 7982
rect 48974 8034 49026 8046
rect 48974 7970 49026 7982
rect 52894 8034 52946 8046
rect 52894 7970 52946 7982
rect 1344 7866 58731 7900
rect 1344 7814 15520 7866
rect 15572 7814 15624 7866
rect 15676 7814 15728 7866
rect 15780 7814 29827 7866
rect 29879 7814 29931 7866
rect 29983 7814 30035 7866
rect 30087 7814 44134 7866
rect 44186 7814 44238 7866
rect 44290 7814 44342 7866
rect 44394 7814 58441 7866
rect 58493 7814 58545 7866
rect 58597 7814 58649 7866
rect 58701 7814 58731 7866
rect 1344 7780 58731 7814
rect 1822 7698 1874 7710
rect 1822 7634 1874 7646
rect 5294 7698 5346 7710
rect 5294 7634 5346 7646
rect 5630 7698 5682 7710
rect 5630 7634 5682 7646
rect 7534 7698 7586 7710
rect 7534 7634 7586 7646
rect 7982 7698 8034 7710
rect 7982 7634 8034 7646
rect 8430 7698 8482 7710
rect 8430 7634 8482 7646
rect 9438 7698 9490 7710
rect 9438 7634 9490 7646
rect 9662 7698 9714 7710
rect 9662 7634 9714 7646
rect 18174 7698 18226 7710
rect 18174 7634 18226 7646
rect 24670 7698 24722 7710
rect 24670 7634 24722 7646
rect 34862 7698 34914 7710
rect 34862 7634 34914 7646
rect 41022 7698 41074 7710
rect 45278 7698 45330 7710
rect 43586 7646 43598 7698
rect 43650 7646 43662 7698
rect 41022 7634 41074 7646
rect 45278 7634 45330 7646
rect 46062 7698 46114 7710
rect 46062 7634 46114 7646
rect 46398 7698 46450 7710
rect 46398 7634 46450 7646
rect 47182 7698 47234 7710
rect 47182 7634 47234 7646
rect 48862 7698 48914 7710
rect 48862 7634 48914 7646
rect 12126 7586 12178 7598
rect 25678 7586 25730 7598
rect 3378 7534 3390 7586
rect 3442 7534 3454 7586
rect 3826 7534 3838 7586
rect 3890 7534 3902 7586
rect 14018 7534 14030 7586
rect 14082 7534 14094 7586
rect 12126 7522 12178 7534
rect 25678 7522 25730 7534
rect 25790 7586 25842 7598
rect 30830 7586 30882 7598
rect 27458 7534 27470 7586
rect 27522 7534 27534 7586
rect 25790 7522 25842 7534
rect 30830 7522 30882 7534
rect 34190 7586 34242 7598
rect 40910 7586 40962 7598
rect 38770 7534 38782 7586
rect 38834 7534 38846 7586
rect 34190 7522 34242 7534
rect 40910 7522 40962 7534
rect 41246 7586 41298 7598
rect 45054 7586 45106 7598
rect 42130 7534 42142 7586
rect 42194 7534 42206 7586
rect 44706 7534 44718 7586
rect 44770 7534 44782 7586
rect 41246 7522 41298 7534
rect 45054 7522 45106 7534
rect 45838 7586 45890 7598
rect 45838 7522 45890 7534
rect 46958 7586 47010 7598
rect 46958 7522 47010 7534
rect 2830 7474 2882 7486
rect 2830 7410 2882 7422
rect 4062 7474 4114 7486
rect 4062 7410 4114 7422
rect 4398 7474 4450 7486
rect 7086 7474 7138 7486
rect 6178 7422 6190 7474
rect 6242 7422 6254 7474
rect 4398 7410 4450 7422
rect 7086 7410 7138 7422
rect 9774 7474 9826 7486
rect 9774 7410 9826 7422
rect 10334 7474 10386 7486
rect 11230 7474 11282 7486
rect 10546 7422 10558 7474
rect 10610 7422 10622 7474
rect 10334 7410 10386 7422
rect 11230 7410 11282 7422
rect 11902 7474 11954 7486
rect 11902 7410 11954 7422
rect 12574 7474 12626 7486
rect 17838 7474 17890 7486
rect 12898 7422 12910 7474
rect 12962 7422 12974 7474
rect 14578 7422 14590 7474
rect 14642 7422 14654 7474
rect 15362 7422 15374 7474
rect 15426 7422 15438 7474
rect 12574 7410 12626 7422
rect 17838 7410 17890 7422
rect 18174 7474 18226 7486
rect 18174 7410 18226 7422
rect 18510 7474 18562 7486
rect 18510 7410 18562 7422
rect 20190 7474 20242 7486
rect 21086 7474 21138 7486
rect 28926 7474 28978 7486
rect 20402 7422 20414 7474
rect 20466 7422 20478 7474
rect 26002 7422 26014 7474
rect 26066 7422 26078 7474
rect 27682 7422 27694 7474
rect 27746 7422 27758 7474
rect 28242 7422 28254 7474
rect 28306 7422 28318 7474
rect 20190 7410 20242 7422
rect 21086 7410 21138 7422
rect 28926 7410 28978 7422
rect 29934 7474 29986 7486
rect 34526 7474 34578 7486
rect 30258 7422 30270 7474
rect 30322 7422 30334 7474
rect 29934 7410 29986 7422
rect 34526 7410 34578 7422
rect 34750 7474 34802 7486
rect 45726 7474 45778 7486
rect 40114 7422 40126 7474
rect 40178 7422 40190 7474
rect 42018 7422 42030 7474
rect 42082 7422 42094 7474
rect 43698 7422 43710 7474
rect 43762 7422 43774 7474
rect 34750 7410 34802 7422
rect 45726 7410 45778 7422
rect 46286 7474 46338 7486
rect 46286 7410 46338 7422
rect 46622 7474 46674 7486
rect 46622 7410 46674 7422
rect 46846 7474 46898 7486
rect 58046 7474 58098 7486
rect 57138 7422 57150 7474
rect 57202 7422 57214 7474
rect 46846 7410 46898 7422
rect 58046 7410 58098 7422
rect 13358 7362 13410 7374
rect 2370 7310 2382 7362
rect 2434 7310 2446 7362
rect 6514 7310 6526 7362
rect 6578 7310 6590 7362
rect 12226 7310 12238 7362
rect 12290 7310 12302 7362
rect 13358 7298 13410 7310
rect 15934 7362 15986 7374
rect 48078 7362 48130 7374
rect 57598 7362 57650 7374
rect 45378 7310 45390 7362
rect 45442 7310 45454 7362
rect 56802 7310 56814 7362
rect 56866 7310 56878 7362
rect 15934 7298 15986 7310
rect 48078 7298 48130 7310
rect 57598 7298 57650 7310
rect 29038 7250 29090 7262
rect 7186 7198 7198 7250
rect 7250 7247 7262 7250
rect 7746 7247 7758 7250
rect 7250 7201 7758 7247
rect 7250 7198 7262 7201
rect 7746 7198 7758 7201
rect 7810 7198 7822 7250
rect 25218 7198 25230 7250
rect 25282 7198 25294 7250
rect 29038 7186 29090 7198
rect 33966 7250 34018 7262
rect 57934 7250 57986 7262
rect 39106 7198 39118 7250
rect 39170 7198 39182 7250
rect 33966 7186 34018 7198
rect 57934 7186 57986 7198
rect 1344 7082 58576 7116
rect 1344 7030 8367 7082
rect 8419 7030 8471 7082
rect 8523 7030 8575 7082
rect 8627 7030 22674 7082
rect 22726 7030 22778 7082
rect 22830 7030 22882 7082
rect 22934 7030 36981 7082
rect 37033 7030 37085 7082
rect 37137 7030 37189 7082
rect 37241 7030 51288 7082
rect 51340 7030 51392 7082
rect 51444 7030 51496 7082
rect 51548 7030 58576 7082
rect 1344 6996 58576 7030
rect 3614 6914 3666 6926
rect 27918 6914 27970 6926
rect 43934 6914 43986 6926
rect 3266 6862 3278 6914
rect 3330 6862 3342 6914
rect 4386 6862 4398 6914
rect 4450 6911 4462 6914
rect 4834 6911 4846 6914
rect 4450 6865 4846 6911
rect 4450 6862 4462 6865
rect 4834 6862 4846 6865
rect 4898 6862 4910 6914
rect 16146 6862 16158 6914
rect 16210 6862 16222 6914
rect 27570 6862 27582 6914
rect 27634 6862 27646 6914
rect 35634 6862 35646 6914
rect 35698 6862 35710 6914
rect 43138 6862 43150 6914
rect 43202 6862 43214 6914
rect 3614 6850 3666 6862
rect 27918 6850 27970 6862
rect 43934 6850 43986 6862
rect 44270 6914 44322 6926
rect 52782 6914 52834 6926
rect 46834 6862 46846 6914
rect 46898 6862 46910 6914
rect 44270 6850 44322 6862
rect 52782 6850 52834 6862
rect 2718 6802 2770 6814
rect 2718 6738 2770 6750
rect 4398 6802 4450 6814
rect 4398 6738 4450 6750
rect 4734 6802 4786 6814
rect 7758 6802 7810 6814
rect 6514 6750 6526 6802
rect 6578 6750 6590 6802
rect 4734 6738 4786 6750
rect 7758 6738 7810 6750
rect 9998 6802 10050 6814
rect 28142 6802 28194 6814
rect 15586 6750 15598 6802
rect 15650 6750 15662 6802
rect 17490 6750 17502 6802
rect 17554 6750 17566 6802
rect 24210 6750 24222 6802
rect 24274 6750 24286 6802
rect 35410 6750 35422 6802
rect 35474 6750 35486 6802
rect 42690 6750 42702 6802
rect 42754 6750 42766 6802
rect 51090 6750 51102 6802
rect 51154 6750 51166 6802
rect 55010 6750 55022 6802
rect 55074 6750 55086 6802
rect 9998 6738 10050 6750
rect 28142 6738 28194 6750
rect 3838 6690 3890 6702
rect 1698 6638 1710 6690
rect 1762 6638 1774 6690
rect 3838 6626 3890 6638
rect 5742 6690 5794 6702
rect 18174 6690 18226 6702
rect 33070 6690 33122 6702
rect 6402 6638 6414 6690
rect 6466 6638 6478 6690
rect 7522 6638 7534 6690
rect 7586 6638 7598 6690
rect 15922 6638 15934 6690
rect 15986 6638 15998 6690
rect 16370 6638 16382 6690
rect 16434 6638 16446 6690
rect 17378 6638 17390 6690
rect 17442 6638 17454 6690
rect 18498 6638 18510 6690
rect 18562 6638 18574 6690
rect 24098 6638 24110 6690
rect 24162 6638 24174 6690
rect 5742 6626 5794 6638
rect 18174 6626 18226 6638
rect 33070 6626 33122 6638
rect 33966 6690 34018 6702
rect 33966 6626 34018 6638
rect 34638 6690 34690 6702
rect 40910 6690 40962 6702
rect 35186 6638 35198 6690
rect 35250 6638 35262 6690
rect 38210 6638 38222 6690
rect 38274 6638 38286 6690
rect 39218 6638 39230 6690
rect 39282 6638 39294 6690
rect 34638 6626 34690 6638
rect 40910 6626 40962 6638
rect 41246 6690 41298 6702
rect 46734 6690 46786 6702
rect 48526 6690 48578 6702
rect 42018 6638 42030 6690
rect 42082 6638 42094 6690
rect 42802 6638 42814 6690
rect 42866 6638 42878 6690
rect 44258 6638 44270 6690
rect 44322 6638 44334 6690
rect 44818 6638 44830 6690
rect 44882 6638 44894 6690
rect 46050 6638 46062 6690
rect 46114 6638 46126 6690
rect 47170 6638 47182 6690
rect 47234 6638 47246 6690
rect 41246 6626 41298 6638
rect 46734 6626 46786 6638
rect 48526 6626 48578 6638
rect 48750 6690 48802 6702
rect 57038 6690 57090 6702
rect 48962 6638 48974 6690
rect 49026 6638 49038 6690
rect 50754 6638 50766 6690
rect 50818 6638 50830 6690
rect 54898 6638 54910 6690
rect 54962 6638 54974 6690
rect 55346 6638 55358 6690
rect 55410 6638 55422 6690
rect 48750 6626 48802 6638
rect 57038 6626 57090 6638
rect 57374 6690 57426 6702
rect 57374 6626 57426 6638
rect 18062 6578 18114 6590
rect 6178 6526 6190 6578
rect 6242 6526 6254 6578
rect 18062 6514 18114 6526
rect 25006 6578 25058 6590
rect 25006 6514 25058 6526
rect 25118 6578 25170 6590
rect 25118 6514 25170 6526
rect 32734 6578 32786 6590
rect 32734 6514 32786 6526
rect 33630 6578 33682 6590
rect 33630 6514 33682 6526
rect 33742 6578 33794 6590
rect 33742 6514 33794 6526
rect 39006 6578 39058 6590
rect 39006 6514 39058 6526
rect 52670 6578 52722 6590
rect 52670 6514 52722 6526
rect 7870 6466 7922 6478
rect 7870 6402 7922 6414
rect 23886 6466 23938 6478
rect 23886 6402 23938 6414
rect 24782 6466 24834 6478
rect 24782 6402 24834 6414
rect 32398 6466 32450 6478
rect 32398 6402 32450 6414
rect 32846 6466 32898 6478
rect 32846 6402 32898 6414
rect 50094 6466 50146 6478
rect 50094 6402 50146 6414
rect 51998 6466 52050 6478
rect 51998 6402 52050 6414
rect 52782 6466 52834 6478
rect 52782 6402 52834 6414
rect 1344 6298 58731 6332
rect 1344 6246 15520 6298
rect 15572 6246 15624 6298
rect 15676 6246 15728 6298
rect 15780 6246 29827 6298
rect 29879 6246 29931 6298
rect 29983 6246 30035 6298
rect 30087 6246 44134 6298
rect 44186 6246 44238 6298
rect 44290 6246 44342 6298
rect 44394 6246 58441 6298
rect 58493 6246 58545 6298
rect 58597 6246 58649 6298
rect 58701 6246 58731 6298
rect 1344 6212 58731 6246
rect 1822 6130 1874 6142
rect 1822 6066 1874 6078
rect 3502 6130 3554 6142
rect 3502 6066 3554 6078
rect 4734 6130 4786 6142
rect 4734 6066 4786 6078
rect 5070 6130 5122 6142
rect 5070 6066 5122 6078
rect 5518 6130 5570 6142
rect 5518 6066 5570 6078
rect 6638 6130 6690 6142
rect 6638 6066 6690 6078
rect 6974 6130 7026 6142
rect 6974 6066 7026 6078
rect 7758 6130 7810 6142
rect 7758 6066 7810 6078
rect 8430 6130 8482 6142
rect 8430 6066 8482 6078
rect 19294 6130 19346 6142
rect 19294 6066 19346 6078
rect 21758 6130 21810 6142
rect 21758 6066 21810 6078
rect 25342 6130 25394 6142
rect 25342 6066 25394 6078
rect 28254 6130 28306 6142
rect 28254 6066 28306 6078
rect 28814 6130 28866 6142
rect 28814 6066 28866 6078
rect 36990 6130 37042 6142
rect 36990 6066 37042 6078
rect 37550 6130 37602 6142
rect 39902 6130 39954 6142
rect 38210 6078 38222 6130
rect 38274 6078 38286 6130
rect 37550 6066 37602 6078
rect 39902 6066 39954 6078
rect 40126 6130 40178 6142
rect 40126 6066 40178 6078
rect 42142 6130 42194 6142
rect 51326 6130 51378 6142
rect 50642 6078 50654 6130
rect 50706 6078 50718 6130
rect 42142 6066 42194 6078
rect 51326 6066 51378 6078
rect 51662 6130 51714 6142
rect 51662 6066 51714 6078
rect 52222 6130 52274 6142
rect 56142 6130 56194 6142
rect 54002 6078 54014 6130
rect 54066 6078 54078 6130
rect 52222 6066 52274 6078
rect 56142 6066 56194 6078
rect 18398 6018 18450 6030
rect 18398 5954 18450 5966
rect 19070 6018 19122 6030
rect 19070 5954 19122 5966
rect 21422 6018 21474 6030
rect 21422 5954 21474 5966
rect 27358 6018 27410 6030
rect 27358 5954 27410 5966
rect 33294 6018 33346 6030
rect 50094 6018 50146 6030
rect 38434 5966 38446 6018
rect 38498 5966 38510 6018
rect 43026 5966 43038 6018
rect 43090 5966 43102 6018
rect 48066 5966 48078 6018
rect 48130 5966 48142 6018
rect 33294 5954 33346 5966
rect 50094 5954 50146 5966
rect 50990 6018 51042 6030
rect 50990 5954 51042 5966
rect 51102 6018 51154 6030
rect 51102 5954 51154 5966
rect 52110 6018 52162 6030
rect 52110 5954 52162 5966
rect 2606 5906 2658 5918
rect 2606 5842 2658 5854
rect 8206 5906 8258 5918
rect 8206 5842 8258 5854
rect 8318 5906 8370 5918
rect 8318 5842 8370 5854
rect 8766 5906 8818 5918
rect 8766 5842 8818 5854
rect 10222 5906 10274 5918
rect 10222 5842 10274 5854
rect 10446 5906 10498 5918
rect 10446 5842 10498 5854
rect 10670 5906 10722 5918
rect 10670 5842 10722 5854
rect 18846 5906 18898 5918
rect 18846 5842 18898 5854
rect 19406 5906 19458 5918
rect 19406 5842 19458 5854
rect 21646 5906 21698 5918
rect 21646 5842 21698 5854
rect 22094 5906 22146 5918
rect 22094 5842 22146 5854
rect 22430 5906 22482 5918
rect 27806 5906 27858 5918
rect 31950 5906 32002 5918
rect 27010 5854 27022 5906
rect 27074 5854 27086 5906
rect 31714 5854 31726 5906
rect 31778 5854 31790 5906
rect 22430 5842 22482 5854
rect 27806 5842 27858 5854
rect 31950 5842 32002 5854
rect 32398 5906 32450 5918
rect 32398 5842 32450 5854
rect 34974 5906 35026 5918
rect 34974 5842 35026 5854
rect 35198 5906 35250 5918
rect 35198 5842 35250 5854
rect 35646 5906 35698 5918
rect 39790 5906 39842 5918
rect 48862 5906 48914 5918
rect 37874 5854 37886 5906
rect 37938 5854 37950 5906
rect 38322 5854 38334 5906
rect 38386 5854 38398 5906
rect 42018 5854 42030 5906
rect 42082 5854 42094 5906
rect 42802 5854 42814 5906
rect 42866 5854 42878 5906
rect 46834 5854 46846 5906
rect 46898 5854 46910 5906
rect 47058 5854 47070 5906
rect 47122 5854 47134 5906
rect 47618 5854 47630 5906
rect 47682 5854 47694 5906
rect 35646 5842 35698 5854
rect 39790 5842 39842 5854
rect 48862 5842 48914 5854
rect 48974 5906 49026 5918
rect 48974 5842 49026 5854
rect 49086 5906 49138 5918
rect 49534 5906 49586 5918
rect 49186 5854 49198 5906
rect 49250 5854 49262 5906
rect 49086 5842 49138 5854
rect 49534 5842 49586 5854
rect 50318 5906 50370 5918
rect 55694 5906 55746 5918
rect 58046 5906 58098 5918
rect 54002 5854 54014 5906
rect 54066 5854 54078 5906
rect 54338 5854 54350 5906
rect 54402 5854 54414 5906
rect 56914 5854 56926 5906
rect 56978 5854 56990 5906
rect 50318 5842 50370 5854
rect 55694 5842 55746 5854
rect 58046 5842 58098 5854
rect 2382 5794 2434 5806
rect 2382 5730 2434 5742
rect 3838 5794 3890 5806
rect 3838 5730 3890 5742
rect 6078 5794 6130 5806
rect 6078 5730 6130 5742
rect 10558 5794 10610 5806
rect 10558 5730 10610 5742
rect 35086 5794 35138 5806
rect 55246 5794 55298 5806
rect 42690 5742 42702 5794
rect 42754 5742 42766 5794
rect 53890 5742 53902 5794
rect 53954 5742 53966 5794
rect 35086 5730 35138 5742
rect 55246 5730 55298 5742
rect 55470 5794 55522 5806
rect 55470 5730 55522 5742
rect 2942 5682 2994 5694
rect 18510 5682 18562 5694
rect 5058 5630 5070 5682
rect 5122 5679 5134 5682
rect 6066 5679 6078 5682
rect 5122 5633 6078 5679
rect 5122 5630 5134 5633
rect 6066 5630 6078 5633
rect 6130 5630 6142 5682
rect 2942 5618 2994 5630
rect 18510 5618 18562 5630
rect 27022 5682 27074 5694
rect 27022 5618 27074 5630
rect 32174 5682 32226 5694
rect 32174 5618 32226 5630
rect 32510 5682 32562 5694
rect 32510 5618 32562 5630
rect 33070 5682 33122 5694
rect 33070 5618 33122 5630
rect 33406 5682 33458 5694
rect 33406 5618 33458 5630
rect 52222 5682 52274 5694
rect 52222 5618 52274 5630
rect 1344 5514 58576 5548
rect 1344 5462 8367 5514
rect 8419 5462 8471 5514
rect 8523 5462 8575 5514
rect 8627 5462 22674 5514
rect 22726 5462 22778 5514
rect 22830 5462 22882 5514
rect 22934 5462 36981 5514
rect 37033 5462 37085 5514
rect 37137 5462 37189 5514
rect 37241 5462 51288 5514
rect 51340 5462 51392 5514
rect 51444 5462 51496 5514
rect 51548 5462 58576 5514
rect 1344 5428 58576 5462
rect 18958 5346 19010 5358
rect 4722 5294 4734 5346
rect 4786 5294 4798 5346
rect 11666 5294 11678 5346
rect 11730 5294 11742 5346
rect 18958 5282 19010 5294
rect 28254 5346 28306 5358
rect 28254 5282 28306 5294
rect 28478 5346 28530 5358
rect 28478 5282 28530 5294
rect 29598 5346 29650 5358
rect 29598 5282 29650 5294
rect 35086 5346 35138 5358
rect 35086 5282 35138 5294
rect 35758 5346 35810 5358
rect 35758 5282 35810 5294
rect 38334 5346 38386 5358
rect 49198 5346 49250 5358
rect 47058 5294 47070 5346
rect 47122 5294 47134 5346
rect 38334 5282 38386 5294
rect 49198 5282 49250 5294
rect 2270 5234 2322 5246
rect 2270 5170 2322 5182
rect 2718 5234 2770 5246
rect 2718 5170 2770 5182
rect 3166 5234 3218 5246
rect 8206 5234 8258 5246
rect 12686 5234 12738 5246
rect 22542 5234 22594 5246
rect 27246 5234 27298 5246
rect 31502 5234 31554 5246
rect 7298 5182 7310 5234
rect 7362 5182 7374 5234
rect 10770 5182 10782 5234
rect 10834 5182 10846 5234
rect 13794 5182 13806 5234
rect 13858 5182 13870 5234
rect 19282 5182 19294 5234
rect 19346 5182 19358 5234
rect 23986 5182 23998 5234
rect 24050 5182 24062 5234
rect 30594 5182 30606 5234
rect 30658 5182 30670 5234
rect 3166 5170 3218 5182
rect 8206 5170 8258 5182
rect 12686 5170 12738 5182
rect 22542 5170 22594 5182
rect 27246 5170 27298 5182
rect 31502 5170 31554 5182
rect 34414 5234 34466 5246
rect 34414 5170 34466 5182
rect 34526 5234 34578 5246
rect 34526 5170 34578 5182
rect 34862 5234 34914 5246
rect 34862 5170 34914 5182
rect 35870 5234 35922 5246
rect 35870 5170 35922 5182
rect 37662 5234 37714 5246
rect 37662 5170 37714 5182
rect 38558 5234 38610 5246
rect 38558 5170 38610 5182
rect 41582 5234 41634 5246
rect 41582 5170 41634 5182
rect 43374 5234 43426 5246
rect 49422 5234 49474 5246
rect 48738 5182 48750 5234
rect 48802 5182 48814 5234
rect 43374 5170 43426 5182
rect 49422 5170 49474 5182
rect 49758 5234 49810 5246
rect 49758 5170 49810 5182
rect 50878 5234 50930 5246
rect 50878 5170 50930 5182
rect 51326 5234 51378 5246
rect 51326 5170 51378 5182
rect 55470 5234 55522 5246
rect 55470 5170 55522 5182
rect 8094 5122 8146 5134
rect 1810 5070 1822 5122
rect 1874 5070 1886 5122
rect 3714 5070 3726 5122
rect 3778 5070 3790 5122
rect 4162 5070 4174 5122
rect 4226 5070 4238 5122
rect 4834 5070 4846 5122
rect 4898 5070 4910 5122
rect 5730 5070 5742 5122
rect 5794 5070 5806 5122
rect 6178 5070 6190 5122
rect 6242 5070 6254 5122
rect 8094 5058 8146 5070
rect 8318 5122 8370 5134
rect 8318 5058 8370 5070
rect 8766 5122 8818 5134
rect 16382 5122 16434 5134
rect 20526 5122 20578 5134
rect 9202 5070 9214 5122
rect 9266 5070 9278 5122
rect 10882 5070 10894 5122
rect 10946 5070 10958 5122
rect 13570 5070 13582 5122
rect 13634 5070 13646 5122
rect 15586 5070 15598 5122
rect 15650 5070 15662 5122
rect 20178 5070 20190 5122
rect 20242 5070 20254 5122
rect 8766 5058 8818 5070
rect 16382 5058 16434 5070
rect 20526 5058 20578 5070
rect 20638 5122 20690 5134
rect 20638 5058 20690 5070
rect 23326 5122 23378 5134
rect 23326 5058 23378 5070
rect 23662 5122 23714 5134
rect 27806 5122 27858 5134
rect 25778 5070 25790 5122
rect 25842 5070 25854 5122
rect 23662 5058 23714 5070
rect 27806 5058 27858 5070
rect 28142 5122 28194 5134
rect 43822 5122 43874 5134
rect 29698 5070 29710 5122
rect 29762 5070 29774 5122
rect 30818 5070 30830 5122
rect 30882 5070 30894 5122
rect 39442 5070 39454 5122
rect 39506 5070 39518 5122
rect 39778 5070 39790 5122
rect 39842 5070 39854 5122
rect 40674 5070 40686 5122
rect 40738 5070 40750 5122
rect 43586 5070 43598 5122
rect 43650 5070 43662 5122
rect 28142 5058 28194 5070
rect 43822 5058 43874 5070
rect 45278 5122 45330 5134
rect 55582 5122 55634 5134
rect 57710 5122 57762 5134
rect 45602 5070 45614 5122
rect 45666 5070 45678 5122
rect 46722 5070 46734 5122
rect 46786 5070 46798 5122
rect 48290 5070 48302 5122
rect 48354 5070 48366 5122
rect 54562 5070 54574 5122
rect 54626 5070 54638 5122
rect 57474 5070 57486 5122
rect 57538 5070 57550 5122
rect 45278 5058 45330 5070
rect 55582 5058 55634 5070
rect 57710 5058 57762 5070
rect 19182 5010 19234 5022
rect 4946 4958 4958 5010
rect 5010 4958 5022 5010
rect 9538 4958 9550 5010
rect 9602 4958 9614 5010
rect 13906 4958 13918 5010
rect 13970 4958 13982 5010
rect 15810 4958 15822 5010
rect 15874 4958 15886 5010
rect 19182 4946 19234 4958
rect 25566 5010 25618 5022
rect 25566 4946 25618 4958
rect 29150 5010 29202 5022
rect 29362 4958 29374 5010
rect 29426 4958 29438 5010
rect 39890 4958 39902 5010
rect 39954 4958 39966 5010
rect 29150 4946 29202 4958
rect 12798 4898 12850 4910
rect 12798 4834 12850 4846
rect 16718 4898 16770 4910
rect 16718 4834 16770 4846
rect 20750 4898 20802 4910
rect 20750 4834 20802 4846
rect 27134 4898 27186 4910
rect 27134 4834 27186 4846
rect 27358 4898 27410 4910
rect 27358 4834 27410 4846
rect 28142 4898 28194 4910
rect 28142 4834 28194 4846
rect 29262 4898 29314 4910
rect 39118 4898 39170 4910
rect 44942 4898 44994 4910
rect 35410 4846 35422 4898
rect 35474 4846 35486 4898
rect 37986 4846 37998 4898
rect 38050 4846 38062 4898
rect 40002 4846 40014 4898
rect 40066 4846 40078 4898
rect 29262 4834 29314 4846
rect 39118 4834 39170 4846
rect 44942 4834 44994 4846
rect 49646 4898 49698 4910
rect 49646 4834 49698 4846
rect 49870 4898 49922 4910
rect 49870 4834 49922 4846
rect 50430 4898 50482 4910
rect 50430 4834 50482 4846
rect 1344 4730 58731 4764
rect 1344 4678 15520 4730
rect 15572 4678 15624 4730
rect 15676 4678 15728 4730
rect 15780 4678 29827 4730
rect 29879 4678 29931 4730
rect 29983 4678 30035 4730
rect 30087 4678 44134 4730
rect 44186 4678 44238 4730
rect 44290 4678 44342 4730
rect 44394 4678 58441 4730
rect 58493 4678 58545 4730
rect 58597 4678 58649 4730
rect 58701 4678 58731 4730
rect 1344 4644 58731 4678
rect 2494 4562 2546 4574
rect 2034 4510 2046 4562
rect 2098 4510 2110 4562
rect 2494 4498 2546 4510
rect 3166 4562 3218 4574
rect 3166 4498 3218 4510
rect 4398 4562 4450 4574
rect 4398 4498 4450 4510
rect 4958 4562 5010 4574
rect 4958 4498 5010 4510
rect 5182 4562 5234 4574
rect 5182 4498 5234 4510
rect 5294 4562 5346 4574
rect 5294 4498 5346 4510
rect 5630 4562 5682 4574
rect 9550 4562 9602 4574
rect 6626 4510 6638 4562
rect 6690 4510 6702 4562
rect 5630 4498 5682 4510
rect 9550 4498 9602 4510
rect 9774 4562 9826 4574
rect 9774 4498 9826 4510
rect 13470 4562 13522 4574
rect 13470 4498 13522 4510
rect 19966 4562 20018 4574
rect 19966 4498 20018 4510
rect 23998 4562 24050 4574
rect 23998 4498 24050 4510
rect 24334 4562 24386 4574
rect 24334 4498 24386 4510
rect 25230 4562 25282 4574
rect 25230 4498 25282 4510
rect 25454 4562 25506 4574
rect 28478 4562 28530 4574
rect 27682 4510 27694 4562
rect 27746 4510 27758 4562
rect 25454 4498 25506 4510
rect 28478 4498 28530 4510
rect 36318 4562 36370 4574
rect 36318 4498 36370 4510
rect 40350 4562 40402 4574
rect 47966 4562 48018 4574
rect 44482 4510 44494 4562
rect 44546 4510 44558 4562
rect 40350 4498 40402 4510
rect 47966 4498 48018 4510
rect 48974 4562 49026 4574
rect 48974 4498 49026 4510
rect 55806 4562 55858 4574
rect 55806 4498 55858 4510
rect 56030 4562 56082 4574
rect 56030 4498 56082 4510
rect 58046 4562 58098 4574
rect 58046 4498 58098 4510
rect 8206 4450 8258 4462
rect 8206 4386 8258 4398
rect 9886 4450 9938 4462
rect 9886 4386 9938 4398
rect 12910 4450 12962 4462
rect 16382 4450 16434 4462
rect 19518 4450 19570 4462
rect 14466 4398 14478 4450
rect 14530 4398 14542 4450
rect 16146 4398 16158 4450
rect 16210 4398 16222 4450
rect 18050 4398 18062 4450
rect 18114 4398 18126 4450
rect 12910 4386 12962 4398
rect 16382 4386 16434 4398
rect 19518 4386 19570 4398
rect 19742 4450 19794 4462
rect 19742 4386 19794 4398
rect 20078 4450 20130 4462
rect 20078 4386 20130 4398
rect 20638 4450 20690 4462
rect 22766 4450 22818 4462
rect 21410 4398 21422 4450
rect 21474 4398 21486 4450
rect 20638 4386 20690 4398
rect 22766 4386 22818 4398
rect 24110 4450 24162 4462
rect 24110 4386 24162 4398
rect 25566 4450 25618 4462
rect 25566 4386 25618 4398
rect 26686 4450 26738 4462
rect 26686 4386 26738 4398
rect 30606 4450 30658 4462
rect 30606 4386 30658 4398
rect 32510 4450 32562 4462
rect 32510 4386 32562 4398
rect 33294 4450 33346 4462
rect 38670 4450 38722 4462
rect 37314 4398 37326 4450
rect 37378 4398 37390 4450
rect 33294 4386 33346 4398
rect 38670 4386 38722 4398
rect 41358 4450 41410 4462
rect 47406 4450 47458 4462
rect 45154 4398 45166 4450
rect 45218 4398 45230 4450
rect 41358 4386 41410 4398
rect 47406 4386 47458 4398
rect 47742 4450 47794 4462
rect 47742 4386 47794 4398
rect 51550 4450 51602 4462
rect 51550 4386 51602 4398
rect 4622 4338 4674 4350
rect 1810 4286 1822 4338
rect 1874 4286 1886 4338
rect 4622 4274 4674 4286
rect 6078 4338 6130 4350
rect 6078 4274 6130 4286
rect 6302 4338 6354 4350
rect 10558 4338 10610 4350
rect 12014 4338 12066 4350
rect 13246 4338 13298 4350
rect 7522 4286 7534 4338
rect 7586 4286 7598 4338
rect 7970 4286 7982 4338
rect 8034 4286 8046 4338
rect 10994 4286 11006 4338
rect 11058 4286 11070 4338
rect 12450 4286 12462 4338
rect 12514 4286 12526 4338
rect 6302 4274 6354 4286
rect 10558 4274 10610 4286
rect 12014 4274 12066 4286
rect 13246 4274 13298 4286
rect 13358 4338 13410 4350
rect 18734 4338 18786 4350
rect 22430 4338 22482 4350
rect 13794 4286 13806 4338
rect 13858 4286 13870 4338
rect 17938 4286 17950 4338
rect 18002 4286 18014 4338
rect 20962 4286 20974 4338
rect 21026 4286 21038 4338
rect 13358 4274 13410 4286
rect 18734 4274 18786 4286
rect 22430 4274 22482 4286
rect 22878 4338 22930 4350
rect 24670 4338 24722 4350
rect 27134 4338 27186 4350
rect 23762 4286 23774 4338
rect 23826 4286 23838 4338
rect 25890 4286 25902 4338
rect 25954 4286 25966 4338
rect 22878 4274 22930 4286
rect 24670 4274 24722 4286
rect 27134 4274 27186 4286
rect 28366 4338 28418 4350
rect 28366 4274 28418 4286
rect 28590 4338 28642 4350
rect 28590 4274 28642 4286
rect 29038 4338 29090 4350
rect 29038 4274 29090 4286
rect 30830 4338 30882 4350
rect 33070 4338 33122 4350
rect 41246 4338 41298 4350
rect 31938 4286 31950 4338
rect 32002 4286 32014 4338
rect 32274 4286 32286 4338
rect 32338 4286 32350 4338
rect 37426 4286 37438 4338
rect 37490 4286 37502 4338
rect 39218 4286 39230 4338
rect 39282 4286 39294 4338
rect 30830 4274 30882 4286
rect 33070 4274 33122 4286
rect 41246 4274 41298 4286
rect 41582 4338 41634 4350
rect 49310 4338 49362 4350
rect 57598 4338 57650 4350
rect 42578 4286 42590 4338
rect 42642 4286 42654 4338
rect 43810 4286 43822 4338
rect 43874 4286 43886 4338
rect 44146 4286 44158 4338
rect 44210 4286 44222 4338
rect 49522 4286 49534 4338
rect 49586 4286 49598 4338
rect 51090 4286 51102 4338
rect 51154 4286 51166 4338
rect 55458 4286 55470 4338
rect 55522 4286 55534 4338
rect 57810 4286 57822 4338
rect 57874 4286 57886 4338
rect 41582 4274 41634 4286
rect 49310 4274 49362 4286
rect 57598 4274 57650 4286
rect 3614 4226 3666 4238
rect 3614 4162 3666 4174
rect 4062 4226 4114 4238
rect 4062 4162 4114 4174
rect 11454 4226 11506 4238
rect 31166 4226 31218 4238
rect 14242 4174 14254 4226
rect 14306 4174 14318 4226
rect 26002 4174 26014 4226
rect 26066 4174 26078 4226
rect 26786 4174 26798 4226
rect 26850 4174 26862 4226
rect 11454 4162 11506 4174
rect 31166 4162 31218 4174
rect 33182 4226 33234 4238
rect 50206 4226 50258 4238
rect 55918 4226 55970 4238
rect 38994 4174 39006 4226
rect 39058 4174 39070 4226
rect 48066 4174 48078 4226
rect 48130 4174 48142 4226
rect 50642 4174 50654 4226
rect 50706 4174 50718 4226
rect 33182 4162 33234 4174
rect 50206 4162 50258 4174
rect 55918 4162 55970 4174
rect 19070 4114 19122 4126
rect 3378 4062 3390 4114
rect 3442 4111 3454 4114
rect 3602 4111 3614 4114
rect 3442 4065 3614 4111
rect 3442 4062 3454 4065
rect 3602 4062 3614 4065
rect 3666 4111 3678 4114
rect 4050 4111 4062 4114
rect 3666 4065 4062 4111
rect 3666 4062 3678 4065
rect 4050 4062 4062 4065
rect 4114 4062 4126 4114
rect 19070 4050 19122 4062
rect 20974 4114 21026 4126
rect 23438 4114 23490 4126
rect 21858 4062 21870 4114
rect 21922 4062 21934 4114
rect 20974 4050 21026 4062
rect 23438 4050 23490 4062
rect 23774 4114 23826 4126
rect 23774 4050 23826 4062
rect 26462 4114 26514 4126
rect 26462 4050 26514 4062
rect 27358 4114 27410 4126
rect 27358 4050 27410 4062
rect 36654 4114 36706 4126
rect 36654 4050 36706 4062
rect 1344 3946 58576 3980
rect 1344 3894 8367 3946
rect 8419 3894 8471 3946
rect 8523 3894 8575 3946
rect 8627 3894 22674 3946
rect 22726 3894 22778 3946
rect 22830 3894 22882 3946
rect 22934 3894 36981 3946
rect 37033 3894 37085 3946
rect 37137 3894 37189 3946
rect 37241 3894 51288 3946
rect 51340 3894 51392 3946
rect 51444 3894 51496 3946
rect 51548 3894 58576 3946
rect 1344 3860 58576 3894
rect 6862 3778 6914 3790
rect 6862 3714 6914 3726
rect 13470 3778 13522 3790
rect 13470 3714 13522 3726
rect 21870 3778 21922 3790
rect 32958 3778 33010 3790
rect 22194 3726 22206 3778
rect 22258 3726 22270 3778
rect 21870 3714 21922 3726
rect 32958 3714 33010 3726
rect 36542 3778 36594 3790
rect 36542 3714 36594 3726
rect 36878 3778 36930 3790
rect 36878 3714 36930 3726
rect 56814 3778 56866 3790
rect 56814 3714 56866 3726
rect 57038 3778 57090 3790
rect 57038 3714 57090 3726
rect 3502 3666 3554 3678
rect 2818 3614 2830 3666
rect 2882 3614 2894 3666
rect 3502 3602 3554 3614
rect 3950 3666 4002 3678
rect 3950 3602 4002 3614
rect 4734 3666 4786 3678
rect 4734 3602 4786 3614
rect 7198 3666 7250 3678
rect 23662 3666 23714 3678
rect 13234 3614 13246 3666
rect 13298 3614 13310 3666
rect 7198 3602 7250 3614
rect 23662 3602 23714 3614
rect 25678 3666 25730 3678
rect 25678 3602 25730 3614
rect 32286 3666 32338 3678
rect 32286 3602 32338 3614
rect 32846 3666 32898 3678
rect 32846 3602 32898 3614
rect 41246 3666 41298 3678
rect 46846 3666 46898 3678
rect 42018 3614 42030 3666
rect 42082 3614 42094 3666
rect 43922 3614 43934 3666
rect 43986 3614 43998 3666
rect 44706 3614 44718 3666
rect 44770 3614 44782 3666
rect 41246 3602 41298 3614
rect 46846 3602 46898 3614
rect 47630 3666 47682 3678
rect 47630 3602 47682 3614
rect 48190 3666 48242 3678
rect 48190 3602 48242 3614
rect 56590 3666 56642 3678
rect 56590 3602 56642 3614
rect 57486 3666 57538 3678
rect 57486 3602 57538 3614
rect 21646 3554 21698 3566
rect 1698 3502 1710 3554
rect 1762 3502 1774 3554
rect 6290 3502 6302 3554
rect 6354 3502 6366 3554
rect 6514 3502 6526 3554
rect 6578 3502 6590 3554
rect 13122 3502 13134 3554
rect 13186 3502 13198 3554
rect 21646 3490 21698 3502
rect 24558 3554 24610 3566
rect 24558 3490 24610 3502
rect 24894 3554 24946 3566
rect 24894 3490 24946 3502
rect 25118 3554 25170 3566
rect 25118 3490 25170 3502
rect 25566 3554 25618 3566
rect 48526 3554 48578 3566
rect 57934 3554 57986 3566
rect 32610 3502 32622 3554
rect 32674 3502 32686 3554
rect 37538 3502 37550 3554
rect 37602 3502 37614 3554
rect 41458 3502 41470 3554
rect 41522 3502 41534 3554
rect 42354 3502 42366 3554
rect 42418 3502 42430 3554
rect 44818 3502 44830 3554
rect 44882 3502 44894 3554
rect 55570 3502 55582 3554
rect 55634 3502 55646 3554
rect 25566 3490 25618 3502
rect 48526 3490 48578 3502
rect 57934 3490 57986 3502
rect 4286 3442 4338 3454
rect 4286 3378 4338 3390
rect 6750 3442 6802 3454
rect 6750 3378 6802 3390
rect 23774 3442 23826 3454
rect 23774 3378 23826 3390
rect 24670 3442 24722 3454
rect 24670 3378 24722 3390
rect 25790 3442 25842 3454
rect 42702 3442 42754 3454
rect 37650 3390 37662 3442
rect 37714 3390 37726 3442
rect 41906 3390 41918 3442
rect 41970 3390 41982 3442
rect 25790 3378 25842 3390
rect 42702 3378 42754 3390
rect 48974 3442 49026 3454
rect 48974 3378 49026 3390
rect 56254 3442 56306 3454
rect 56254 3378 56306 3390
rect 57598 3442 57650 3454
rect 57598 3378 57650 3390
rect 57822 3442 57874 3454
rect 57822 3378 57874 3390
rect 1344 3162 58731 3196
rect 1344 3110 15520 3162
rect 15572 3110 15624 3162
rect 15676 3110 15728 3162
rect 15780 3110 29827 3162
rect 29879 3110 29931 3162
rect 29983 3110 30035 3162
rect 30087 3110 44134 3162
rect 44186 3110 44238 3162
rect 44290 3110 44342 3162
rect 44394 3110 58441 3162
rect 58493 3110 58545 3162
rect 58597 3110 58649 3162
rect 58701 3110 58731 3162
rect 1344 3076 58731 3110
<< via1 >>
rect 48750 26798 48802 26850
rect 49086 26798 49138 26850
rect 49758 26798 49810 26850
rect 15520 26630 15572 26682
rect 15624 26630 15676 26682
rect 15728 26630 15780 26682
rect 29827 26630 29879 26682
rect 29931 26630 29983 26682
rect 30035 26630 30087 26682
rect 44134 26630 44186 26682
rect 44238 26630 44290 26682
rect 44342 26630 44394 26682
rect 58441 26630 58493 26682
rect 58545 26630 58597 26682
rect 58649 26630 58701 26682
rect 12462 26462 12514 26514
rect 21310 26462 21362 26514
rect 48750 26462 48802 26514
rect 50318 26462 50370 26514
rect 52222 26462 52274 26514
rect 57710 26462 57762 26514
rect 7982 26350 8034 26402
rect 8206 26350 8258 26402
rect 9326 26350 9378 26402
rect 14030 26350 14082 26402
rect 16046 26350 16098 26402
rect 16382 26350 16434 26402
rect 20750 26350 20802 26402
rect 26686 26350 26738 26402
rect 28926 26350 28978 26402
rect 37438 26350 37490 26402
rect 40126 26350 40178 26402
rect 49758 26350 49810 26402
rect 50654 26350 50706 26402
rect 2158 26238 2210 26290
rect 5518 26238 5570 26290
rect 6862 26238 6914 26290
rect 7198 26238 7250 26290
rect 7310 26238 7362 26290
rect 7646 26238 7698 26290
rect 11118 26238 11170 26290
rect 11342 26238 11394 26290
rect 12350 26238 12402 26290
rect 13246 26238 13298 26290
rect 13582 26238 13634 26290
rect 16270 26238 16322 26290
rect 17502 26238 17554 26290
rect 19182 26238 19234 26290
rect 22094 26238 22146 26290
rect 22654 26238 22706 26290
rect 26910 26238 26962 26290
rect 27358 26238 27410 26290
rect 28702 26238 28754 26290
rect 29486 26238 29538 26290
rect 31278 26238 31330 26290
rect 33070 26238 33122 26290
rect 33742 26238 33794 26290
rect 34190 26238 34242 26290
rect 36206 26238 36258 26290
rect 37998 26238 38050 26290
rect 41358 26238 41410 26290
rect 48638 26238 48690 26290
rect 49534 26238 49586 26290
rect 49982 26238 50034 26290
rect 51326 26238 51378 26290
rect 56926 26238 56978 26290
rect 5070 26126 5122 26178
rect 5966 26126 6018 26178
rect 8878 26126 8930 26178
rect 9886 26126 9938 26178
rect 10558 26126 10610 26178
rect 19630 26126 19682 26178
rect 20078 26126 20130 26178
rect 21982 26126 22034 26178
rect 23102 26126 23154 26178
rect 23438 26126 23490 26178
rect 24670 26126 24722 26178
rect 25454 26126 25506 26178
rect 26014 26126 26066 26178
rect 26462 26126 26514 26178
rect 27134 26126 27186 26178
rect 27694 26126 27746 26178
rect 29934 26126 29986 26178
rect 32286 26126 32338 26178
rect 33518 26126 33570 26178
rect 35422 26126 35474 26178
rect 38558 26126 38610 26178
rect 39902 26126 39954 26178
rect 46846 26126 46898 26178
rect 47630 26126 47682 26178
rect 48078 26126 48130 26178
rect 51774 26126 51826 26178
rect 53006 26126 53058 26178
rect 53230 26126 53282 26178
rect 56590 26126 56642 26178
rect 4062 26014 4114 26066
rect 15038 26014 15090 26066
rect 19070 26014 19122 26066
rect 20974 26014 21026 26066
rect 23662 26014 23714 26066
rect 23998 26014 24050 26066
rect 29822 26014 29874 26066
rect 31166 26014 31218 26066
rect 36318 26014 36370 26066
rect 42702 26014 42754 26066
rect 49198 26014 49250 26066
rect 51214 26014 51266 26066
rect 53454 26014 53506 26066
rect 53678 26014 53730 26066
rect 54126 26014 54178 26066
rect 8367 25846 8419 25898
rect 8471 25846 8523 25898
rect 8575 25846 8627 25898
rect 22674 25846 22726 25898
rect 22778 25846 22830 25898
rect 22882 25846 22934 25898
rect 36981 25846 37033 25898
rect 37085 25846 37137 25898
rect 37189 25846 37241 25898
rect 51288 25846 51340 25898
rect 51392 25846 51444 25898
rect 51496 25846 51548 25898
rect 25230 25678 25282 25730
rect 37550 25678 37602 25730
rect 54910 25678 54962 25730
rect 3054 25566 3106 25618
rect 5854 25566 5906 25618
rect 9774 25566 9826 25618
rect 12014 25566 12066 25618
rect 29374 25566 29426 25618
rect 30046 25566 30098 25618
rect 32062 25566 32114 25618
rect 35534 25566 35586 25618
rect 42142 25566 42194 25618
rect 50430 25566 50482 25618
rect 53566 25566 53618 25618
rect 1710 25454 1762 25506
rect 6974 25454 7026 25506
rect 7198 25454 7250 25506
rect 7758 25454 7810 25506
rect 9438 25454 9490 25506
rect 11454 25454 11506 25506
rect 13470 25454 13522 25506
rect 14366 25454 14418 25506
rect 15150 25454 15202 25506
rect 17166 25454 17218 25506
rect 17614 25454 17666 25506
rect 19742 25454 19794 25506
rect 21534 25454 21586 25506
rect 23102 25454 23154 25506
rect 24670 25454 24722 25506
rect 26126 25454 26178 25506
rect 27694 25454 27746 25506
rect 30158 25454 30210 25506
rect 32398 25454 32450 25506
rect 32846 25454 32898 25506
rect 34526 25454 34578 25506
rect 36094 25454 36146 25506
rect 36430 25454 36482 25506
rect 36990 25454 37042 25506
rect 37214 25454 37266 25506
rect 38782 25454 38834 25506
rect 39006 25454 39058 25506
rect 41806 25454 41858 25506
rect 45390 25454 45442 25506
rect 46510 25454 46562 25506
rect 48638 25454 48690 25506
rect 51886 25454 51938 25506
rect 52110 25454 52162 25506
rect 53454 25454 53506 25506
rect 55470 25454 55522 25506
rect 8094 25342 8146 25394
rect 9102 25342 9154 25394
rect 12910 25342 12962 25394
rect 16718 25342 16770 25394
rect 20190 25342 20242 25394
rect 21310 25342 21362 25394
rect 23886 25342 23938 25394
rect 24446 25342 24498 25394
rect 25566 25342 25618 25394
rect 26686 25342 26738 25394
rect 28478 25342 28530 25394
rect 32734 25342 32786 25394
rect 35870 25342 35922 25394
rect 42702 25342 42754 25394
rect 45166 25342 45218 25394
rect 49198 25342 49250 25394
rect 5182 25230 5234 25282
rect 6302 25230 6354 25282
rect 6638 25230 6690 25282
rect 12350 25230 12402 25282
rect 13582 25230 13634 25282
rect 16494 25230 16546 25282
rect 16606 25230 16658 25282
rect 20638 25230 20690 25282
rect 23326 25230 23378 25282
rect 34974 25230 35026 25282
rect 36318 25230 36370 25282
rect 43262 25230 43314 25282
rect 48190 25230 48242 25282
rect 50206 25230 50258 25282
rect 51550 25230 51602 25282
rect 52894 25230 52946 25282
rect 15520 25062 15572 25114
rect 15624 25062 15676 25114
rect 15728 25062 15780 25114
rect 29827 25062 29879 25114
rect 29931 25062 29983 25114
rect 30035 25062 30087 25114
rect 44134 25062 44186 25114
rect 44238 25062 44290 25114
rect 44342 25062 44394 25114
rect 58441 25062 58493 25114
rect 58545 25062 58597 25114
rect 58649 25062 58701 25114
rect 9774 24894 9826 24946
rect 25566 24894 25618 24946
rect 31390 24894 31442 24946
rect 31726 24894 31778 24946
rect 34078 24894 34130 24946
rect 35870 24894 35922 24946
rect 39678 24894 39730 24946
rect 47854 24894 47906 24946
rect 49198 24894 49250 24946
rect 5630 24782 5682 24834
rect 8766 24782 8818 24834
rect 11902 24782 11954 24834
rect 12910 24782 12962 24834
rect 21422 24782 21474 24834
rect 22654 24782 22706 24834
rect 24670 24782 24722 24834
rect 27246 24782 27298 24834
rect 29150 24782 29202 24834
rect 32174 24782 32226 24834
rect 33182 24782 33234 24834
rect 33406 24782 33458 24834
rect 33742 24782 33794 24834
rect 33854 24782 33906 24834
rect 34974 24782 35026 24834
rect 37438 24782 37490 24834
rect 44718 24782 44770 24834
rect 49646 24782 49698 24834
rect 53006 24782 53058 24834
rect 54910 24782 54962 24834
rect 2494 24670 2546 24722
rect 3166 24670 3218 24722
rect 3726 24670 3778 24722
rect 4958 24670 5010 24722
rect 5406 24670 5458 24722
rect 6414 24670 6466 24722
rect 7646 24670 7698 24722
rect 10222 24670 10274 24722
rect 13358 24670 13410 24722
rect 14030 24670 14082 24722
rect 14926 24670 14978 24722
rect 15150 24670 15202 24722
rect 17502 24670 17554 24722
rect 18398 24670 18450 24722
rect 19070 24670 19122 24722
rect 20414 24670 20466 24722
rect 22542 24670 22594 24722
rect 25678 24670 25730 24722
rect 26686 24670 26738 24722
rect 28366 24670 28418 24722
rect 30158 24670 30210 24722
rect 30494 24670 30546 24722
rect 32062 24670 32114 24722
rect 36430 24670 36482 24722
rect 38558 24670 38610 24722
rect 39566 24670 39618 24722
rect 42030 24670 42082 24722
rect 42366 24670 42418 24722
rect 42702 24670 42754 24722
rect 43038 24670 43090 24722
rect 43262 24670 43314 24722
rect 45950 24670 46002 24722
rect 49086 24670 49138 24722
rect 50878 24670 50930 24722
rect 52446 24670 52498 24722
rect 54574 24670 54626 24722
rect 7198 24558 7250 24610
rect 8990 24558 9042 24610
rect 9886 24558 9938 24610
rect 10446 24558 10498 24610
rect 13918 24558 13970 24610
rect 14590 24558 14642 24610
rect 16158 24558 16210 24610
rect 18286 24558 18338 24610
rect 21198 24558 21250 24610
rect 22318 24558 22370 24610
rect 25790 24558 25842 24610
rect 27806 24558 27858 24610
rect 30942 24558 30994 24610
rect 33070 24558 33122 24610
rect 39342 24558 39394 24610
rect 42254 24558 42306 24610
rect 42926 24558 42978 24610
rect 44494 24558 44546 24610
rect 48190 24558 48242 24610
rect 52110 24558 52162 24610
rect 53454 24558 53506 24610
rect 55246 24558 55298 24610
rect 56590 24558 56642 24610
rect 1710 24446 1762 24498
rect 6638 24446 6690 24498
rect 17502 24446 17554 24498
rect 22206 24446 22258 24498
rect 32174 24446 32226 24498
rect 47294 24446 47346 24498
rect 47518 24446 47570 24498
rect 48078 24446 48130 24498
rect 56814 24446 56866 24498
rect 57150 24446 57202 24498
rect 8367 24278 8419 24330
rect 8471 24278 8523 24330
rect 8575 24278 8627 24330
rect 22674 24278 22726 24330
rect 22778 24278 22830 24330
rect 22882 24278 22934 24330
rect 36981 24278 37033 24330
rect 37085 24278 37137 24330
rect 37189 24278 37241 24330
rect 51288 24278 51340 24330
rect 51392 24278 51444 24330
rect 51496 24278 51548 24330
rect 21646 24110 21698 24162
rect 36094 24110 36146 24162
rect 3278 23998 3330 24050
rect 8878 23998 8930 24050
rect 12910 23998 12962 24050
rect 15262 23998 15314 24050
rect 20078 23998 20130 24050
rect 22094 23998 22146 24050
rect 30606 23998 30658 24050
rect 33630 23998 33682 24050
rect 34750 23998 34802 24050
rect 35310 23998 35362 24050
rect 35982 23998 36034 24050
rect 42926 23998 42978 24050
rect 51102 23998 51154 24050
rect 3054 23886 3106 23938
rect 7758 23886 7810 23938
rect 10334 23886 10386 23938
rect 10782 23886 10834 23938
rect 11006 23886 11058 23938
rect 11342 23886 11394 23938
rect 12238 23886 12290 23938
rect 14926 23886 14978 23938
rect 15710 23886 15762 23938
rect 16158 23886 16210 23938
rect 16718 23886 16770 23938
rect 18510 23886 18562 23938
rect 19966 23886 20018 23938
rect 21870 23886 21922 23938
rect 24334 23886 24386 23938
rect 24782 23886 24834 23938
rect 27358 23886 27410 23938
rect 27806 23886 27858 23938
rect 28478 23886 28530 23938
rect 29150 23886 29202 23938
rect 31054 23886 31106 23938
rect 32846 23886 32898 23938
rect 35758 23886 35810 23938
rect 37886 23886 37938 23938
rect 39230 23886 39282 23938
rect 41022 23886 41074 23938
rect 42814 23886 42866 23938
rect 46846 23886 46898 23938
rect 47182 23886 47234 23938
rect 49534 23886 49586 23938
rect 51550 23886 51602 23938
rect 53118 23886 53170 23938
rect 53566 23886 53618 23938
rect 55582 23886 55634 23938
rect 56590 23886 56642 23938
rect 57934 23886 57986 23938
rect 4622 23774 4674 23826
rect 5742 23774 5794 23826
rect 8094 23774 8146 23826
rect 9102 23774 9154 23826
rect 12350 23774 12402 23826
rect 18174 23774 18226 23826
rect 20526 23774 20578 23826
rect 20638 23774 20690 23826
rect 22206 23774 22258 23826
rect 22430 23774 22482 23826
rect 22766 23774 22818 23826
rect 25342 23774 25394 23826
rect 27918 23774 27970 23826
rect 29262 23774 29314 23826
rect 31726 23774 31778 23826
rect 32734 23774 32786 23826
rect 35086 23774 35138 23826
rect 37550 23774 37602 23826
rect 41694 23774 41746 23826
rect 44270 23774 44322 23826
rect 47070 23774 47122 23826
rect 48638 23774 48690 23826
rect 49646 23774 49698 23826
rect 51326 23774 51378 23826
rect 54238 23774 54290 23826
rect 55806 23774 55858 23826
rect 2270 23662 2322 23714
rect 5070 23662 5122 23714
rect 6638 23662 6690 23714
rect 8318 23662 8370 23714
rect 12014 23662 12066 23714
rect 13582 23662 13634 23714
rect 20862 23662 20914 23714
rect 26462 23662 26514 23714
rect 29710 23662 29762 23714
rect 35310 23662 35362 23714
rect 38558 23662 38610 23714
rect 46286 23662 46338 23714
rect 52110 23662 52162 23714
rect 54798 23662 54850 23714
rect 56478 23662 56530 23714
rect 57598 23662 57650 23714
rect 15520 23494 15572 23546
rect 15624 23494 15676 23546
rect 15728 23494 15780 23546
rect 29827 23494 29879 23546
rect 29931 23494 29983 23546
rect 30035 23494 30087 23546
rect 44134 23494 44186 23546
rect 44238 23494 44290 23546
rect 44342 23494 44394 23546
rect 58441 23494 58493 23546
rect 58545 23494 58597 23546
rect 58649 23494 58701 23546
rect 16942 23326 16994 23378
rect 22318 23326 22370 23378
rect 22542 23326 22594 23378
rect 24558 23326 24610 23378
rect 52670 23326 52722 23378
rect 1710 23214 1762 23266
rect 2942 23214 2994 23266
rect 10670 23214 10722 23266
rect 13470 23214 13522 23266
rect 16158 23214 16210 23266
rect 24446 23214 24498 23266
rect 28030 23214 28082 23266
rect 28702 23214 28754 23266
rect 35310 23214 35362 23266
rect 38222 23214 38274 23266
rect 47294 23214 47346 23266
rect 49534 23214 49586 23266
rect 50542 23214 50594 23266
rect 52110 23214 52162 23266
rect 52446 23214 52498 23266
rect 55470 23214 55522 23266
rect 2494 23102 2546 23154
rect 3726 23102 3778 23154
rect 5966 23102 6018 23154
rect 6750 23102 6802 23154
rect 8766 23102 8818 23154
rect 9774 23102 9826 23154
rect 11454 23102 11506 23154
rect 12686 23102 12738 23154
rect 14478 23102 14530 23154
rect 16494 23102 16546 23154
rect 18286 23102 18338 23154
rect 19966 23102 20018 23154
rect 21982 23102 22034 23154
rect 22654 23102 22706 23154
rect 23326 23102 23378 23154
rect 23886 23102 23938 23154
rect 24782 23102 24834 23154
rect 25230 23102 25282 23154
rect 27134 23102 27186 23154
rect 30382 23102 30434 23154
rect 30830 23102 30882 23154
rect 31054 23102 31106 23154
rect 32062 23102 32114 23154
rect 33742 23102 33794 23154
rect 35422 23102 35474 23154
rect 36878 23102 36930 23154
rect 37102 23102 37154 23154
rect 40350 23102 40402 23154
rect 41246 23102 41298 23154
rect 41582 23102 41634 23154
rect 42254 23102 42306 23154
rect 42926 23102 42978 23154
rect 46510 23102 46562 23154
rect 47070 23102 47122 23154
rect 48750 23102 48802 23154
rect 51886 23102 51938 23154
rect 52334 23102 52386 23154
rect 53454 23102 53506 23154
rect 53678 23102 53730 23154
rect 54126 23102 54178 23154
rect 54798 23102 54850 23154
rect 56926 23102 56978 23154
rect 2718 22990 2770 23042
rect 3614 22990 3666 23042
rect 6302 22990 6354 23042
rect 8094 22990 8146 23042
rect 11678 22990 11730 23042
rect 17614 22990 17666 23042
rect 17838 22990 17890 23042
rect 19742 22990 19794 23042
rect 21086 22990 21138 23042
rect 23438 22990 23490 23042
rect 25678 22990 25730 23042
rect 26462 22990 26514 23042
rect 26798 22990 26850 23042
rect 30494 22990 30546 23042
rect 33630 22990 33682 23042
rect 34750 22990 34802 23042
rect 36318 22990 36370 23042
rect 37662 22990 37714 23042
rect 39902 22990 39954 23042
rect 41358 22990 41410 23042
rect 43038 22990 43090 23042
rect 44606 22990 44658 23042
rect 46958 22990 47010 23042
rect 53006 22990 53058 23042
rect 53566 22990 53618 23042
rect 54686 22990 54738 23042
rect 55918 22990 55970 23042
rect 57038 22990 57090 23042
rect 1822 22878 1874 22930
rect 4846 22878 4898 22930
rect 31278 22878 31330 22930
rect 35982 22878 36034 22930
rect 37214 22878 37266 22930
rect 39006 22878 39058 22930
rect 57262 22878 57314 22930
rect 8367 22710 8419 22762
rect 8471 22710 8523 22762
rect 8575 22710 8627 22762
rect 22674 22710 22726 22762
rect 22778 22710 22830 22762
rect 22882 22710 22934 22762
rect 36981 22710 37033 22762
rect 37085 22710 37137 22762
rect 37189 22710 37241 22762
rect 51288 22710 51340 22762
rect 51392 22710 51444 22762
rect 51496 22710 51548 22762
rect 11902 22542 11954 22594
rect 24670 22542 24722 22594
rect 27134 22542 27186 22594
rect 35198 22542 35250 22594
rect 49422 22542 49474 22594
rect 51662 22542 51714 22594
rect 10782 22430 10834 22482
rect 20190 22430 20242 22482
rect 22206 22430 22258 22482
rect 38110 22430 38162 22482
rect 40350 22430 40402 22482
rect 41470 22430 41522 22482
rect 44270 22430 44322 22482
rect 2382 22318 2434 22370
rect 4398 22318 4450 22370
rect 7198 22318 7250 22370
rect 7758 22318 7810 22370
rect 8542 22318 8594 22370
rect 8878 22318 8930 22370
rect 9102 22318 9154 22370
rect 10894 22318 10946 22370
rect 13582 22318 13634 22370
rect 15262 22318 15314 22370
rect 17278 22318 17330 22370
rect 17838 22318 17890 22370
rect 18622 22318 18674 22370
rect 20414 22318 20466 22370
rect 21534 22318 21586 22370
rect 22990 22318 23042 22370
rect 24334 22318 24386 22370
rect 26574 22318 26626 22370
rect 27134 22318 27186 22370
rect 29598 22318 29650 22370
rect 30158 22318 30210 22370
rect 32062 22318 32114 22370
rect 32734 22318 32786 22370
rect 33518 22318 33570 22370
rect 38222 22318 38274 22370
rect 40014 22318 40066 22370
rect 41022 22318 41074 22370
rect 43598 22318 43650 22370
rect 45950 22318 46002 22370
rect 47070 22318 47122 22370
rect 48414 22318 48466 22370
rect 49534 22318 49586 22370
rect 50654 22318 50706 22370
rect 51438 22318 51490 22370
rect 52782 22318 52834 22370
rect 53006 22318 53058 22370
rect 54350 22318 54402 22370
rect 56366 22318 56418 22370
rect 2718 22206 2770 22258
rect 4622 22206 4674 22258
rect 6190 22206 6242 22258
rect 8206 22206 8258 22258
rect 13694 22206 13746 22258
rect 14254 22206 14306 22258
rect 15934 22206 15986 22258
rect 20750 22206 20802 22258
rect 22430 22206 22482 22258
rect 23550 22206 23602 22258
rect 23998 22206 24050 22258
rect 25678 22206 25730 22258
rect 26238 22206 26290 22258
rect 26798 22206 26850 22258
rect 28254 22206 28306 22258
rect 30830 22206 30882 22258
rect 33406 22206 33458 22258
rect 34414 22206 34466 22258
rect 34862 22206 34914 22258
rect 44046 22206 44098 22258
rect 46062 22206 46114 22258
rect 47966 22206 48018 22258
rect 53230 22206 53282 22258
rect 53678 22206 53730 22258
rect 53790 22206 53842 22258
rect 55470 22206 55522 22258
rect 57486 22206 57538 22258
rect 3390 22094 3442 22146
rect 8318 22094 8370 22146
rect 13022 22094 13074 22146
rect 13806 22094 13858 22146
rect 15038 22094 15090 22146
rect 22766 22094 22818 22146
rect 25342 22094 25394 22146
rect 35534 22094 35586 22146
rect 46958 22094 47010 22146
rect 51998 22094 52050 22146
rect 52894 22094 52946 22146
rect 54014 22094 54066 22146
rect 56478 22094 56530 22146
rect 15520 21926 15572 21978
rect 15624 21926 15676 21978
rect 15728 21926 15780 21978
rect 29827 21926 29879 21978
rect 29931 21926 29983 21978
rect 30035 21926 30087 21978
rect 44134 21926 44186 21978
rect 44238 21926 44290 21978
rect 44342 21926 44394 21978
rect 58441 21926 58493 21978
rect 58545 21926 58597 21978
rect 58649 21926 58701 21978
rect 3390 21758 3442 21810
rect 8878 21758 8930 21810
rect 12798 21758 12850 21810
rect 17726 21758 17778 21810
rect 22766 21758 22818 21810
rect 26574 21758 26626 21810
rect 52334 21758 52386 21810
rect 54238 21758 54290 21810
rect 6974 21646 7026 21698
rect 7422 21646 7474 21698
rect 7982 21646 8034 21698
rect 11902 21646 11954 21698
rect 14366 21646 14418 21698
rect 19630 21646 19682 21698
rect 23662 21646 23714 21698
rect 24558 21646 24610 21698
rect 26462 21646 26514 21698
rect 28590 21646 28642 21698
rect 31390 21646 31442 21698
rect 36990 21646 37042 21698
rect 42142 21646 42194 21698
rect 45278 21646 45330 21698
rect 47406 21646 47458 21698
rect 49310 21646 49362 21698
rect 51438 21646 51490 21698
rect 53902 21646 53954 21698
rect 54462 21646 54514 21698
rect 56030 21646 56082 21698
rect 57710 21646 57762 21698
rect 1710 21534 1762 21586
rect 3502 21534 3554 21586
rect 3838 21534 3890 21586
rect 6078 21534 6130 21586
rect 7198 21534 7250 21586
rect 8318 21534 8370 21586
rect 8990 21534 9042 21586
rect 10222 21534 10274 21586
rect 10670 21534 10722 21586
rect 11790 21534 11842 21586
rect 13918 21534 13970 21586
rect 16046 21534 16098 21586
rect 16270 21534 16322 21586
rect 17614 21534 17666 21586
rect 17950 21534 18002 21586
rect 19854 21534 19906 21586
rect 20414 21534 20466 21586
rect 20862 21534 20914 21586
rect 23102 21534 23154 21586
rect 23886 21534 23938 21586
rect 25230 21534 25282 21586
rect 27694 21534 27746 21586
rect 28702 21534 28754 21586
rect 29710 21534 29762 21586
rect 31054 21534 31106 21586
rect 31838 21534 31890 21586
rect 32286 21534 32338 21586
rect 34414 21534 34466 21586
rect 35870 21534 35922 21586
rect 37550 21534 37602 21586
rect 38334 21534 38386 21586
rect 38782 21534 38834 21586
rect 42030 21534 42082 21586
rect 42366 21534 42418 21586
rect 44046 21534 44098 21586
rect 44718 21534 44770 21586
rect 46622 21534 46674 21586
rect 47182 21534 47234 21586
rect 48750 21534 48802 21586
rect 48974 21534 49026 21586
rect 50990 21534 51042 21586
rect 53342 21534 53394 21586
rect 53790 21534 53842 21586
rect 55246 21534 55298 21586
rect 55470 21534 55522 21586
rect 55806 21534 55858 21586
rect 57262 21534 57314 21586
rect 57934 21534 57986 21586
rect 2718 21422 2770 21474
rect 5966 21422 6018 21474
rect 10334 21422 10386 21474
rect 11454 21422 11506 21474
rect 24334 21422 24386 21474
rect 25678 21422 25730 21474
rect 30158 21422 30210 21474
rect 31950 21422 32002 21474
rect 40238 21422 40290 21474
rect 41134 21422 41186 21474
rect 41470 21422 41522 21474
rect 43710 21422 43762 21474
rect 47630 21422 47682 21474
rect 48190 21422 48242 21474
rect 50654 21422 50706 21474
rect 52782 21422 52834 21474
rect 56702 21422 56754 21474
rect 58046 21422 58098 21474
rect 3390 21310 3442 21362
rect 6414 21310 6466 21362
rect 10110 21310 10162 21362
rect 16046 21310 16098 21362
rect 21422 21310 21474 21362
rect 24670 21310 24722 21362
rect 36766 21310 36818 21362
rect 45054 21310 45106 21362
rect 55694 21310 55746 21362
rect 8367 21142 8419 21194
rect 8471 21142 8523 21194
rect 8575 21142 8627 21194
rect 22674 21142 22726 21194
rect 22778 21142 22830 21194
rect 22882 21142 22934 21194
rect 36981 21142 37033 21194
rect 37085 21142 37137 21194
rect 37189 21142 37241 21194
rect 51288 21142 51340 21194
rect 51392 21142 51444 21194
rect 51496 21142 51548 21194
rect 4958 20974 5010 21026
rect 23662 20974 23714 21026
rect 34862 20974 34914 21026
rect 42142 20974 42194 21026
rect 54350 20974 54402 21026
rect 55246 20974 55298 21026
rect 6302 20862 6354 20914
rect 18510 20862 18562 20914
rect 27022 20862 27074 20914
rect 34526 20862 34578 20914
rect 36430 20862 36482 20914
rect 38558 20862 38610 20914
rect 48078 20862 48130 20914
rect 52894 20862 52946 20914
rect 53790 20862 53842 20914
rect 54798 20862 54850 20914
rect 56478 20862 56530 20914
rect 1822 20750 1874 20802
rect 2606 20750 2658 20802
rect 4734 20750 4786 20802
rect 6750 20750 6802 20802
rect 8430 20750 8482 20802
rect 9662 20750 9714 20802
rect 11566 20750 11618 20802
rect 12798 20750 12850 20802
rect 14030 20750 14082 20802
rect 16046 20750 16098 20802
rect 17054 20750 17106 20802
rect 20414 20750 20466 20802
rect 20638 20750 20690 20802
rect 20750 20750 20802 20802
rect 21534 20750 21586 20802
rect 23326 20750 23378 20802
rect 23998 20750 24050 20802
rect 25118 20750 25170 20802
rect 28254 20750 28306 20802
rect 29150 20750 29202 20802
rect 30382 20750 30434 20802
rect 31838 20750 31890 20802
rect 32174 20750 32226 20802
rect 32398 20750 32450 20802
rect 37214 20750 37266 20802
rect 38782 20750 38834 20802
rect 41134 20750 41186 20802
rect 41918 20750 41970 20802
rect 42702 20750 42754 20802
rect 42814 20750 42866 20802
rect 45838 20750 45890 20802
rect 46062 20750 46114 20802
rect 46734 20750 46786 20802
rect 47406 20750 47458 20802
rect 48526 20750 48578 20802
rect 49534 20750 49586 20802
rect 51550 20750 51602 20802
rect 52670 20750 52722 20802
rect 53118 20750 53170 20802
rect 54014 20750 54066 20802
rect 55022 20750 55074 20802
rect 55694 20750 55746 20802
rect 57710 20750 57762 20802
rect 57934 20750 57986 20802
rect 58158 20750 58210 20802
rect 2942 20638 2994 20690
rect 3278 20638 3330 20690
rect 4622 20638 4674 20690
rect 6862 20638 6914 20690
rect 11006 20638 11058 20690
rect 14590 20638 14642 20690
rect 16606 20638 16658 20690
rect 22542 20638 22594 20690
rect 25006 20638 25058 20690
rect 26574 20638 26626 20690
rect 28366 20638 28418 20690
rect 29374 20638 29426 20690
rect 29822 20638 29874 20690
rect 30494 20638 30546 20690
rect 34190 20638 34242 20690
rect 35086 20638 35138 20690
rect 36990 20638 37042 20690
rect 40350 20638 40402 20690
rect 44046 20638 44098 20690
rect 46958 20638 47010 20690
rect 48862 20638 48914 20690
rect 49198 20638 49250 20690
rect 50878 20638 50930 20690
rect 51886 20638 51938 20690
rect 52222 20638 52274 20690
rect 56814 20638 56866 20690
rect 2270 20526 2322 20578
rect 5854 20526 5906 20578
rect 7758 20526 7810 20578
rect 12798 20526 12850 20578
rect 15038 20526 15090 20578
rect 22654 20526 22706 20578
rect 30718 20526 30770 20578
rect 31054 20526 31106 20578
rect 32846 20526 32898 20578
rect 34414 20526 34466 20578
rect 34974 20526 35026 20578
rect 51998 20526 52050 20578
rect 53230 20526 53282 20578
rect 53342 20526 53394 20578
rect 57374 20526 57426 20578
rect 15520 20358 15572 20410
rect 15624 20358 15676 20410
rect 15728 20358 15780 20410
rect 29827 20358 29879 20410
rect 29931 20358 29983 20410
rect 30035 20358 30087 20410
rect 44134 20358 44186 20410
rect 44238 20358 44290 20410
rect 44342 20358 44394 20410
rect 58441 20358 58493 20410
rect 58545 20358 58597 20410
rect 58649 20358 58701 20410
rect 16830 20190 16882 20242
rect 22766 20190 22818 20242
rect 55918 20190 55970 20242
rect 2158 20078 2210 20130
rect 4622 20078 4674 20130
rect 9774 20078 9826 20130
rect 9998 20078 10050 20130
rect 10334 20078 10386 20130
rect 16270 20078 16322 20130
rect 21870 20078 21922 20130
rect 23326 20078 23378 20130
rect 24222 20078 24274 20130
rect 30494 20078 30546 20130
rect 30606 20078 30658 20130
rect 36318 20078 36370 20130
rect 43822 20078 43874 20130
rect 44158 20078 44210 20130
rect 45054 20078 45106 20130
rect 47070 20078 47122 20130
rect 47518 20078 47570 20130
rect 49198 20078 49250 20130
rect 50094 20078 50146 20130
rect 54014 20078 54066 20130
rect 57710 20078 57762 20130
rect 2046 19966 2098 20018
rect 2942 19966 2994 20018
rect 3166 19966 3218 20018
rect 5182 19966 5234 20018
rect 7758 19966 7810 20018
rect 10558 19966 10610 20018
rect 12574 19966 12626 20018
rect 12910 19966 12962 20018
rect 14814 19966 14866 20018
rect 15598 19966 15650 20018
rect 17390 19966 17442 20018
rect 21310 19966 21362 20018
rect 24446 19966 24498 20018
rect 25566 19966 25618 20018
rect 25902 19966 25954 20018
rect 27470 19966 27522 20018
rect 28590 19966 28642 20018
rect 30046 19966 30098 20018
rect 33070 19966 33122 20018
rect 34190 19966 34242 20018
rect 35310 19966 35362 20018
rect 36094 19966 36146 20018
rect 37886 19966 37938 20018
rect 39678 19966 39730 20018
rect 40238 19966 40290 20018
rect 42030 19966 42082 20018
rect 42366 19966 42418 20018
rect 44494 19966 44546 20018
rect 46286 19966 46338 20018
rect 47742 19966 47794 20018
rect 49422 19966 49474 20018
rect 50878 19966 50930 20018
rect 51102 19966 51154 20018
rect 52894 19966 52946 20018
rect 53566 19966 53618 20018
rect 53902 19966 53954 20018
rect 55134 19966 55186 20018
rect 55246 19966 55298 20018
rect 55470 19966 55522 20018
rect 56926 19966 56978 20018
rect 4846 19854 4898 19906
rect 7086 19854 7138 19906
rect 7646 19854 7698 19906
rect 8878 19854 8930 19906
rect 9886 19854 9938 19906
rect 15822 19854 15874 19906
rect 16494 19854 16546 19906
rect 19518 19854 19570 19906
rect 21086 19854 21138 19906
rect 37326 19854 37378 19906
rect 38894 19854 38946 19906
rect 39342 19854 39394 19906
rect 41470 19854 41522 19906
rect 43262 19854 43314 19906
rect 48974 19854 49026 19906
rect 49310 19854 49362 19906
rect 2046 19742 2098 19794
rect 10782 19742 10834 19794
rect 23662 19742 23714 19794
rect 29486 19742 29538 19794
rect 30494 19742 30546 19794
rect 35646 19742 35698 19794
rect 46174 19742 46226 19794
rect 48078 19742 48130 19794
rect 48750 19742 48802 19794
rect 8367 19574 8419 19626
rect 8471 19574 8523 19626
rect 8575 19574 8627 19626
rect 22674 19574 22726 19626
rect 22778 19574 22830 19626
rect 22882 19574 22934 19626
rect 36981 19574 37033 19626
rect 37085 19574 37137 19626
rect 37189 19574 37241 19626
rect 51288 19574 51340 19626
rect 51392 19574 51444 19626
rect 51496 19574 51548 19626
rect 11006 19406 11058 19458
rect 15038 19406 15090 19458
rect 23774 19406 23826 19458
rect 26238 19406 26290 19458
rect 35198 19406 35250 19458
rect 36206 19406 36258 19458
rect 43934 19406 43986 19458
rect 45054 19406 45106 19458
rect 45950 19406 46002 19458
rect 53454 19406 53506 19458
rect 15598 19294 15650 19346
rect 16942 19294 16994 19346
rect 19406 19294 19458 19346
rect 21422 19294 21474 19346
rect 25118 19294 25170 19346
rect 25902 19294 25954 19346
rect 27022 19294 27074 19346
rect 30270 19294 30322 19346
rect 32398 19294 32450 19346
rect 37550 19294 37602 19346
rect 40574 19294 40626 19346
rect 49646 19294 49698 19346
rect 51662 19294 51714 19346
rect 53118 19294 53170 19346
rect 1710 19182 1762 19234
rect 3614 19182 3666 19234
rect 3950 19182 4002 19234
rect 5742 19182 5794 19234
rect 5854 19182 5906 19234
rect 9326 19182 9378 19234
rect 10110 19182 10162 19234
rect 11230 19182 11282 19234
rect 14254 19182 14306 19234
rect 15710 19182 15762 19234
rect 17054 19182 17106 19234
rect 17614 19182 17666 19234
rect 21534 19182 21586 19234
rect 23326 19182 23378 19234
rect 23998 19182 24050 19234
rect 25006 19182 25058 19234
rect 25566 19182 25618 19234
rect 27694 19182 27746 19234
rect 29150 19182 29202 19234
rect 29374 19182 29426 19234
rect 31166 19182 31218 19234
rect 32622 19182 32674 19234
rect 33518 19182 33570 19234
rect 34078 19182 34130 19234
rect 35870 19182 35922 19234
rect 37102 19182 37154 19234
rect 39006 19182 39058 19234
rect 41134 19182 41186 19234
rect 41806 19182 41858 19234
rect 43150 19182 43202 19234
rect 46062 19182 46114 19234
rect 47294 19182 47346 19234
rect 47966 19182 48018 19234
rect 49198 19182 49250 19234
rect 49870 19182 49922 19234
rect 50878 19182 50930 19234
rect 53230 19182 53282 19234
rect 53342 19182 53394 19234
rect 54350 19182 54402 19234
rect 58158 19182 58210 19234
rect 2270 19070 2322 19122
rect 4622 19070 4674 19122
rect 7646 19070 7698 19122
rect 8542 19070 8594 19122
rect 8766 19070 8818 19122
rect 10558 19070 10610 19122
rect 11454 19070 11506 19122
rect 16494 19070 16546 19122
rect 18174 19070 18226 19122
rect 23214 19070 23266 19122
rect 24558 19070 24610 19122
rect 26014 19070 26066 19122
rect 28030 19070 28082 19122
rect 33854 19070 33906 19122
rect 36094 19070 36146 19122
rect 37214 19070 37266 19122
rect 40462 19070 40514 19122
rect 43038 19070 43090 19122
rect 45278 19070 45330 19122
rect 49198 19070 49250 19122
rect 49422 19070 49474 19122
rect 54462 19070 54514 19122
rect 56254 19070 56306 19122
rect 57598 19070 57650 19122
rect 5070 18958 5122 19010
rect 9102 18958 9154 19010
rect 19630 18958 19682 19010
rect 20638 18958 20690 19010
rect 22766 18958 22818 19010
rect 24110 18958 24162 19010
rect 45166 18958 45218 19010
rect 49758 18958 49810 19010
rect 15520 18790 15572 18842
rect 15624 18790 15676 18842
rect 15728 18790 15780 18842
rect 29827 18790 29879 18842
rect 29931 18790 29983 18842
rect 30035 18790 30087 18842
rect 44134 18790 44186 18842
rect 44238 18790 44290 18842
rect 44342 18790 44394 18842
rect 58441 18790 58493 18842
rect 58545 18790 58597 18842
rect 58649 18790 58701 18842
rect 2158 18622 2210 18674
rect 4398 18622 4450 18674
rect 14814 18622 14866 18674
rect 26350 18622 26402 18674
rect 26910 18622 26962 18674
rect 28702 18622 28754 18674
rect 35086 18622 35138 18674
rect 35870 18622 35922 18674
rect 39230 18622 39282 18674
rect 41470 18622 41522 18674
rect 41694 18622 41746 18674
rect 45166 18622 45218 18674
rect 51886 18622 51938 18674
rect 3614 18510 3666 18562
rect 3950 18510 4002 18562
rect 5742 18510 5794 18562
rect 6750 18510 6802 18562
rect 14702 18510 14754 18562
rect 18846 18510 18898 18562
rect 19742 18510 19794 18562
rect 23102 18510 23154 18562
rect 25566 18510 25618 18562
rect 26462 18510 26514 18562
rect 28030 18510 28082 18562
rect 34974 18510 35026 18562
rect 35758 18510 35810 18562
rect 37102 18510 37154 18562
rect 41246 18510 41298 18562
rect 44718 18510 44770 18562
rect 48862 18510 48914 18562
rect 52334 18510 52386 18562
rect 54462 18510 54514 18562
rect 2046 18398 2098 18450
rect 2830 18398 2882 18450
rect 3838 18398 3890 18450
rect 4174 18398 4226 18450
rect 4510 18398 4562 18450
rect 5294 18398 5346 18450
rect 6078 18398 6130 18450
rect 6974 18398 7026 18450
rect 8654 18398 8706 18450
rect 9886 18398 9938 18450
rect 10222 18398 10274 18450
rect 11566 18398 11618 18450
rect 11902 18398 11954 18450
rect 13694 18398 13746 18450
rect 15822 18398 15874 18450
rect 17390 18398 17442 18450
rect 18398 18398 18450 18450
rect 20750 18398 20802 18450
rect 22542 18398 22594 18450
rect 25230 18398 25282 18450
rect 26126 18398 26178 18450
rect 27358 18398 27410 18450
rect 29150 18398 29202 18450
rect 29598 18398 29650 18450
rect 30494 18398 30546 18450
rect 30830 18398 30882 18450
rect 33182 18398 33234 18450
rect 33406 18398 33458 18450
rect 33854 18398 33906 18450
rect 36094 18398 36146 18450
rect 36318 18398 36370 18450
rect 36654 18398 36706 18450
rect 37214 18398 37266 18450
rect 38782 18398 38834 18450
rect 42814 18398 42866 18450
rect 42926 18398 42978 18450
rect 43598 18398 43650 18450
rect 45502 18398 45554 18450
rect 46398 18398 46450 18450
rect 46734 18398 46786 18450
rect 47070 18398 47122 18450
rect 49198 18398 49250 18450
rect 50542 18398 50594 18450
rect 52558 18398 52610 18450
rect 53902 18398 53954 18450
rect 54798 18398 54850 18450
rect 54910 18398 54962 18450
rect 2494 18286 2546 18338
rect 6302 18286 6354 18338
rect 8990 18286 9042 18338
rect 9662 18286 9714 18338
rect 11230 18286 11282 18338
rect 18062 18286 18114 18338
rect 20974 18286 21026 18338
rect 21534 18286 21586 18338
rect 22318 18286 22370 18338
rect 24670 18286 24722 18338
rect 25902 18286 25954 18338
rect 30718 18286 30770 18338
rect 34526 18286 34578 18338
rect 36542 18286 36594 18338
rect 40350 18286 40402 18338
rect 41358 18286 41410 18338
rect 42142 18286 42194 18338
rect 55806 18286 55858 18338
rect 7982 18174 8034 18226
rect 10670 18174 10722 18226
rect 16158 18174 16210 18226
rect 22206 18174 22258 18226
rect 31166 18174 31218 18226
rect 33070 18174 33122 18226
rect 33630 18174 33682 18226
rect 35198 18174 35250 18226
rect 42254 18174 42306 18226
rect 8367 18006 8419 18058
rect 8471 18006 8523 18058
rect 8575 18006 8627 18058
rect 22674 18006 22726 18058
rect 22778 18006 22830 18058
rect 22882 18006 22934 18058
rect 36981 18006 37033 18058
rect 37085 18006 37137 18058
rect 37189 18006 37241 18058
rect 51288 18006 51340 18058
rect 51392 18006 51444 18058
rect 51496 18006 51548 18058
rect 19518 17838 19570 17890
rect 28478 17838 28530 17890
rect 32622 17838 32674 17890
rect 42254 17838 42306 17890
rect 43262 17838 43314 17890
rect 2942 17726 2994 17778
rect 3726 17726 3778 17778
rect 4286 17726 4338 17778
rect 6078 17726 6130 17778
rect 7198 17726 7250 17778
rect 11006 17726 11058 17778
rect 12014 17726 12066 17778
rect 15038 17726 15090 17778
rect 17390 17726 17442 17778
rect 20190 17726 20242 17778
rect 39118 17726 39170 17778
rect 40910 17726 40962 17778
rect 41806 17726 41858 17778
rect 42590 17726 42642 17778
rect 45278 17726 45330 17778
rect 45614 17726 45666 17778
rect 53118 17726 53170 17778
rect 57374 17726 57426 17778
rect 1822 17614 1874 17666
rect 2270 17614 2322 17666
rect 6862 17614 6914 17666
rect 7086 17614 7138 17666
rect 7982 17614 8034 17666
rect 8206 17614 8258 17666
rect 8318 17614 8370 17666
rect 10222 17614 10274 17666
rect 10446 17614 10498 17666
rect 12350 17614 12402 17666
rect 12910 17614 12962 17666
rect 14030 17614 14082 17666
rect 15150 17614 15202 17666
rect 17502 17614 17554 17666
rect 18174 17614 18226 17666
rect 19294 17614 19346 17666
rect 20302 17614 20354 17666
rect 23438 17614 23490 17666
rect 23774 17614 23826 17666
rect 26238 17614 26290 17666
rect 28366 17614 28418 17666
rect 31502 17614 31554 17666
rect 32174 17614 32226 17666
rect 33294 17614 33346 17666
rect 37550 17614 37602 17666
rect 37774 17614 37826 17666
rect 39790 17614 39842 17666
rect 41470 17614 41522 17666
rect 41694 17614 41746 17666
rect 41918 17614 41970 17666
rect 45054 17614 45106 17666
rect 46286 17614 46338 17666
rect 47630 17614 47682 17666
rect 48302 17614 48354 17666
rect 50878 17614 50930 17666
rect 52782 17614 52834 17666
rect 53342 17614 53394 17666
rect 54238 17614 54290 17666
rect 54574 17614 54626 17666
rect 55694 17614 55746 17666
rect 3390 17502 3442 17554
rect 3614 17502 3666 17554
rect 5742 17502 5794 17554
rect 5966 17502 6018 17554
rect 9662 17502 9714 17554
rect 15822 17502 15874 17554
rect 20526 17502 20578 17554
rect 21758 17502 21810 17554
rect 24334 17502 24386 17554
rect 27694 17502 27746 17554
rect 37102 17502 37154 17554
rect 41246 17502 41298 17554
rect 43038 17502 43090 17554
rect 49422 17502 49474 17554
rect 49758 17502 49810 17554
rect 52894 17502 52946 17554
rect 53566 17502 53618 17554
rect 55134 17502 55186 17554
rect 56142 17502 56194 17554
rect 4734 17390 4786 17442
rect 25342 17390 25394 17442
rect 42478 17390 42530 17442
rect 43150 17390 43202 17442
rect 51214 17390 51266 17442
rect 51662 17390 51714 17442
rect 55022 17390 55074 17442
rect 57038 17390 57090 17442
rect 15520 17222 15572 17274
rect 15624 17222 15676 17274
rect 15728 17222 15780 17274
rect 29827 17222 29879 17274
rect 29931 17222 29983 17274
rect 30035 17222 30087 17274
rect 44134 17222 44186 17274
rect 44238 17222 44290 17274
rect 44342 17222 44394 17274
rect 58441 17222 58493 17274
rect 58545 17222 58597 17274
rect 58649 17222 58701 17274
rect 12686 17054 12738 17106
rect 27918 17054 27970 17106
rect 35758 17054 35810 17106
rect 40238 17054 40290 17106
rect 40462 17054 40514 17106
rect 41022 17054 41074 17106
rect 42142 17054 42194 17106
rect 45390 17054 45442 17106
rect 48078 17054 48130 17106
rect 48862 17054 48914 17106
rect 49310 17054 49362 17106
rect 53454 17054 53506 17106
rect 55470 17054 55522 17106
rect 8430 16942 8482 16994
rect 9550 16942 9602 16994
rect 11006 16942 11058 16994
rect 12014 16942 12066 16994
rect 15598 16942 15650 16994
rect 22766 16942 22818 16994
rect 23326 16942 23378 16994
rect 26462 16942 26514 16994
rect 30718 16942 30770 16994
rect 33070 16942 33122 16994
rect 34302 16942 34354 16994
rect 35198 16942 35250 16994
rect 36206 16942 36258 16994
rect 37550 16942 37602 16994
rect 43598 16942 43650 16994
rect 44270 16942 44322 16994
rect 47182 16942 47234 16994
rect 47518 16942 47570 16994
rect 50990 16942 51042 16994
rect 51886 16942 51938 16994
rect 53902 16942 53954 16994
rect 55918 16942 55970 16994
rect 57710 16942 57762 16994
rect 4174 16830 4226 16882
rect 5630 16830 5682 16882
rect 6526 16830 6578 16882
rect 7086 16830 7138 16882
rect 8878 16830 8930 16882
rect 9662 16830 9714 16882
rect 12686 16830 12738 16882
rect 14590 16830 14642 16882
rect 15038 16830 15090 16882
rect 17390 16830 17442 16882
rect 17614 16830 17666 16882
rect 19294 16830 19346 16882
rect 20414 16830 20466 16882
rect 22542 16830 22594 16882
rect 23550 16830 23602 16882
rect 23998 16830 24050 16882
rect 26014 16830 26066 16882
rect 26238 16830 26290 16882
rect 26350 16830 26402 16882
rect 27358 16830 27410 16882
rect 27694 16830 27746 16882
rect 28366 16830 28418 16882
rect 29262 16830 29314 16882
rect 29598 16830 29650 16882
rect 31054 16830 31106 16882
rect 32062 16830 32114 16882
rect 33294 16830 33346 16882
rect 34638 16830 34690 16882
rect 34974 16830 35026 16882
rect 36094 16830 36146 16882
rect 37102 16830 37154 16882
rect 38894 16830 38946 16882
rect 40126 16830 40178 16882
rect 41134 16830 41186 16882
rect 42478 16830 42530 16882
rect 43486 16830 43538 16882
rect 44606 16830 44658 16882
rect 51326 16830 51378 16882
rect 53342 16830 53394 16882
rect 55694 16830 55746 16882
rect 57038 16830 57090 16882
rect 57934 16830 57986 16882
rect 58158 16830 58210 16882
rect 2046 16718 2098 16770
rect 5518 16718 5570 16770
rect 8094 16718 8146 16770
rect 19742 16718 19794 16770
rect 22430 16718 22482 16770
rect 27246 16718 27298 16770
rect 27806 16718 27858 16770
rect 31726 16718 31778 16770
rect 35086 16718 35138 16770
rect 36766 16718 36818 16770
rect 39230 16718 39282 16770
rect 39454 16718 39506 16770
rect 41246 16718 41298 16770
rect 44158 16718 44210 16770
rect 47742 16718 47794 16770
rect 56926 16718 56978 16770
rect 2270 16606 2322 16658
rect 2494 16606 2546 16658
rect 2718 16606 2770 16658
rect 3166 16606 3218 16658
rect 4734 16606 4786 16658
rect 16606 16606 16658 16658
rect 24334 16606 24386 16658
rect 26910 16606 26962 16658
rect 27022 16606 27074 16658
rect 31278 16606 31330 16658
rect 33518 16606 33570 16658
rect 33742 16606 33794 16658
rect 37774 16606 37826 16658
rect 38110 16606 38162 16658
rect 55358 16606 55410 16658
rect 57262 16606 57314 16658
rect 57598 16606 57650 16658
rect 8367 16438 8419 16490
rect 8471 16438 8523 16490
rect 8575 16438 8627 16490
rect 22674 16438 22726 16490
rect 22778 16438 22830 16490
rect 22882 16438 22934 16490
rect 36981 16438 37033 16490
rect 37085 16438 37137 16490
rect 37189 16438 37241 16490
rect 51288 16438 51340 16490
rect 51392 16438 51444 16490
rect 51496 16438 51548 16490
rect 3390 16270 3442 16322
rect 4398 16270 4450 16322
rect 21310 16270 21362 16322
rect 21646 16270 21698 16322
rect 23438 16270 23490 16322
rect 31166 16270 31218 16322
rect 54014 16270 54066 16322
rect 56142 16270 56194 16322
rect 6078 16158 6130 16210
rect 7982 16158 8034 16210
rect 9998 16158 10050 16210
rect 10894 16158 10946 16210
rect 17726 16158 17778 16210
rect 31390 16158 31442 16210
rect 36430 16158 36482 16210
rect 37774 16158 37826 16210
rect 40462 16158 40514 16210
rect 41694 16158 41746 16210
rect 45166 16158 45218 16210
rect 51438 16158 51490 16210
rect 54574 16158 54626 16210
rect 55582 16158 55634 16210
rect 2270 16046 2322 16098
rect 3054 16046 3106 16098
rect 6526 16046 6578 16098
rect 7086 16046 7138 16098
rect 8542 16046 8594 16098
rect 9662 16046 9714 16098
rect 12350 16046 12402 16098
rect 13470 16046 13522 16098
rect 15262 16046 15314 16098
rect 17950 16046 18002 16098
rect 18734 16046 18786 16098
rect 20078 16046 20130 16098
rect 22206 16046 22258 16098
rect 22766 16046 22818 16098
rect 23214 16046 23266 16098
rect 24558 16046 24610 16098
rect 26126 16046 26178 16098
rect 26574 16046 26626 16098
rect 27134 16046 27186 16098
rect 27918 16046 27970 16098
rect 28366 16046 28418 16098
rect 30046 16046 30098 16098
rect 30382 16046 30434 16098
rect 36990 16046 37042 16098
rect 37662 16046 37714 16098
rect 38782 16046 38834 16098
rect 43710 16046 43762 16098
rect 43934 16046 43986 16098
rect 44382 16046 44434 16098
rect 45054 16046 45106 16098
rect 47630 16046 47682 16098
rect 47854 16046 47906 16098
rect 48974 16046 49026 16098
rect 49310 16046 49362 16098
rect 51102 16046 51154 16098
rect 52110 16046 52162 16098
rect 53678 16046 53730 16098
rect 54910 16046 54962 16098
rect 55806 16046 55858 16098
rect 57374 16046 57426 16098
rect 4622 15934 4674 15986
rect 11230 15934 11282 15986
rect 12686 15934 12738 15986
rect 14478 15934 14530 15986
rect 16606 15934 16658 15986
rect 17166 15934 17218 15986
rect 21534 15934 21586 15986
rect 21982 15934 22034 15986
rect 24334 15934 24386 15986
rect 27358 15934 27410 15986
rect 30158 15934 30210 15986
rect 34862 15934 34914 15986
rect 35086 15934 35138 15986
rect 38222 15934 38274 15986
rect 39230 15934 39282 15986
rect 46510 15934 46562 15986
rect 48078 15934 48130 15986
rect 53230 15934 53282 15986
rect 53454 15934 53506 15986
rect 55022 15934 55074 15986
rect 1710 15822 1762 15874
rect 4510 15822 4562 15874
rect 15038 15822 15090 15874
rect 16270 15822 16322 15874
rect 16494 15822 16546 15874
rect 26686 15822 26738 15874
rect 26910 15822 26962 15874
rect 28478 15822 28530 15874
rect 30830 15822 30882 15874
rect 34974 15822 35026 15874
rect 40238 15822 40290 15874
rect 43822 15822 43874 15874
rect 55246 15822 55298 15874
rect 15520 15654 15572 15706
rect 15624 15654 15676 15706
rect 15728 15654 15780 15706
rect 29827 15654 29879 15706
rect 29931 15654 29983 15706
rect 30035 15654 30087 15706
rect 44134 15654 44186 15706
rect 44238 15654 44290 15706
rect 44342 15654 44394 15706
rect 58441 15654 58493 15706
rect 58545 15654 58597 15706
rect 58649 15654 58701 15706
rect 6750 15486 6802 15538
rect 7422 15486 7474 15538
rect 7870 15486 7922 15538
rect 8878 15486 8930 15538
rect 10110 15486 10162 15538
rect 11566 15486 11618 15538
rect 18734 15486 18786 15538
rect 23102 15486 23154 15538
rect 23326 15486 23378 15538
rect 24446 15486 24498 15538
rect 27918 15486 27970 15538
rect 28142 15486 28194 15538
rect 28254 15486 28306 15538
rect 37102 15486 37154 15538
rect 39006 15486 39058 15538
rect 42142 15486 42194 15538
rect 42590 15486 42642 15538
rect 44606 15486 44658 15538
rect 44830 15486 44882 15538
rect 45390 15486 45442 15538
rect 45838 15486 45890 15538
rect 48078 15486 48130 15538
rect 52110 15486 52162 15538
rect 55246 15486 55298 15538
rect 2606 15374 2658 15426
rect 4398 15374 4450 15426
rect 5294 15374 5346 15426
rect 6638 15374 6690 15426
rect 9662 15374 9714 15426
rect 10558 15374 10610 15426
rect 15486 15374 15538 15426
rect 16046 15374 16098 15426
rect 18062 15374 18114 15426
rect 22318 15374 22370 15426
rect 23886 15374 23938 15426
rect 27022 15374 27074 15426
rect 27694 15374 27746 15426
rect 38110 15374 38162 15426
rect 41694 15374 41746 15426
rect 45726 15374 45778 15426
rect 47854 15374 47906 15426
rect 50654 15374 50706 15426
rect 50990 15374 51042 15426
rect 54686 15374 54738 15426
rect 58046 15374 58098 15426
rect 2382 15262 2434 15314
rect 3054 15262 3106 15314
rect 6078 15262 6130 15314
rect 6974 15262 7026 15314
rect 8990 15262 9042 15314
rect 9550 15262 9602 15314
rect 10670 15262 10722 15314
rect 11454 15262 11506 15314
rect 12350 15262 12402 15314
rect 13918 15262 13970 15314
rect 14142 15262 14194 15314
rect 16270 15262 16322 15314
rect 16382 15262 16434 15314
rect 17726 15262 17778 15314
rect 18622 15262 18674 15314
rect 19182 15262 19234 15314
rect 19518 15262 19570 15314
rect 21534 15262 21586 15314
rect 23438 15262 23490 15314
rect 25230 15262 25282 15314
rect 25454 15262 25506 15314
rect 30830 15262 30882 15314
rect 31054 15262 31106 15314
rect 32062 15262 32114 15314
rect 32510 15262 32562 15314
rect 33966 15262 34018 15314
rect 34190 15262 34242 15314
rect 34414 15262 34466 15314
rect 34638 15262 34690 15314
rect 34974 15262 35026 15314
rect 35198 15262 35250 15314
rect 36990 15262 37042 15314
rect 37886 15262 37938 15314
rect 41134 15262 41186 15314
rect 42366 15262 42418 15314
rect 44270 15262 44322 15314
rect 47518 15262 47570 15314
rect 48974 15262 49026 15314
rect 49198 15262 49250 15314
rect 51214 15262 51266 15314
rect 51438 15262 51490 15314
rect 51662 15262 51714 15314
rect 53454 15262 53506 15314
rect 53678 15262 53730 15314
rect 54126 15262 54178 15314
rect 57150 15262 57202 15314
rect 2046 15150 2098 15202
rect 14254 15150 14306 15202
rect 22094 15150 22146 15202
rect 24110 15150 24162 15202
rect 28254 15150 28306 15202
rect 31726 15150 31778 15202
rect 33518 15150 33570 15202
rect 38334 15150 38386 15202
rect 39342 15150 39394 15202
rect 41582 15150 41634 15202
rect 42478 15150 42530 15202
rect 48190 15150 48242 15202
rect 48750 15150 48802 15202
rect 53902 15150 53954 15202
rect 55806 15150 55858 15202
rect 6078 15038 6130 15090
rect 7086 15038 7138 15090
rect 7422 15038 7474 15090
rect 7646 15038 7698 15090
rect 7982 15038 8034 15090
rect 35646 15038 35698 15090
rect 44494 15038 44546 15090
rect 45838 15038 45890 15090
rect 8367 14870 8419 14922
rect 8471 14870 8523 14922
rect 8575 14870 8627 14922
rect 22674 14870 22726 14922
rect 22778 14870 22830 14922
rect 22882 14870 22934 14922
rect 36981 14870 37033 14922
rect 37085 14870 37137 14922
rect 37189 14870 37241 14922
rect 51288 14870 51340 14922
rect 51392 14870 51444 14922
rect 51496 14870 51548 14922
rect 8654 14702 8706 14754
rect 8990 14702 9042 14754
rect 24222 14702 24274 14754
rect 28366 14702 28418 14754
rect 33518 14702 33570 14754
rect 38670 14702 38722 14754
rect 6302 14590 6354 14642
rect 7646 14590 7698 14642
rect 8430 14590 8482 14642
rect 12126 14590 12178 14642
rect 13582 14590 13634 14642
rect 18734 14590 18786 14642
rect 21870 14590 21922 14642
rect 22430 14590 22482 14642
rect 23662 14590 23714 14642
rect 23886 14590 23938 14642
rect 33070 14590 33122 14642
rect 34750 14590 34802 14642
rect 37886 14590 37938 14642
rect 39566 14590 39618 14642
rect 41470 14590 41522 14642
rect 53454 14590 53506 14642
rect 2606 14478 2658 14530
rect 2942 14478 2994 14530
rect 3950 14478 4002 14530
rect 4286 14478 4338 14530
rect 7534 14478 7586 14530
rect 10782 14478 10834 14530
rect 11006 14478 11058 14530
rect 11342 14478 11394 14530
rect 11566 14478 11618 14530
rect 12238 14478 12290 14530
rect 16046 14478 16098 14530
rect 18174 14478 18226 14530
rect 18622 14478 18674 14530
rect 21646 14478 21698 14530
rect 22654 14478 22706 14530
rect 22878 14478 22930 14530
rect 24446 14478 24498 14530
rect 24782 14478 24834 14530
rect 27470 14478 27522 14530
rect 30718 14478 30770 14530
rect 31166 14478 31218 14530
rect 32958 14478 33010 14530
rect 34862 14478 34914 14530
rect 35758 14478 35810 14530
rect 37998 14478 38050 14530
rect 38222 14478 38274 14530
rect 40574 14478 40626 14530
rect 41358 14478 41410 14530
rect 41694 14478 41746 14530
rect 44830 14478 44882 14530
rect 45054 14478 45106 14530
rect 48190 14478 48242 14530
rect 49198 14478 49250 14530
rect 50878 14478 50930 14530
rect 51214 14478 51266 14530
rect 51438 14478 51490 14530
rect 53006 14478 53058 14530
rect 53230 14478 53282 14530
rect 54462 14478 54514 14530
rect 56478 14478 56530 14530
rect 2270 14366 2322 14418
rect 4398 14366 4450 14418
rect 4734 14366 4786 14418
rect 8094 14366 8146 14418
rect 9550 14366 9602 14418
rect 12910 14366 12962 14418
rect 14254 14366 14306 14418
rect 14590 14366 14642 14418
rect 16382 14366 16434 14418
rect 17166 14366 17218 14418
rect 19742 14366 19794 14418
rect 23214 14366 23266 14418
rect 26014 14366 26066 14418
rect 27134 14366 27186 14418
rect 28366 14366 28418 14418
rect 28478 14366 28530 14418
rect 35870 14366 35922 14418
rect 39230 14366 39282 14418
rect 45278 14366 45330 14418
rect 47518 14366 47570 14418
rect 49086 14366 49138 14418
rect 55022 14366 55074 14418
rect 57038 14366 57090 14418
rect 1710 14254 1762 14306
rect 2718 14254 2770 14306
rect 4846 14254 4898 14306
rect 5070 14254 5122 14306
rect 5854 14254 5906 14306
rect 9214 14254 9266 14306
rect 9438 14254 9490 14306
rect 10446 14254 10498 14306
rect 11118 14254 11170 14306
rect 23102 14254 23154 14306
rect 26798 14254 26850 14306
rect 27246 14254 27298 14306
rect 27806 14254 27858 14306
rect 34750 14254 34802 14306
rect 36094 14254 36146 14306
rect 39454 14254 39506 14306
rect 40686 14254 40738 14306
rect 40910 14254 40962 14306
rect 41918 14254 41970 14306
rect 44942 14254 44994 14306
rect 48526 14254 48578 14306
rect 49982 14254 50034 14306
rect 50542 14254 50594 14306
rect 51102 14254 51154 14306
rect 52110 14254 52162 14306
rect 52558 14254 52610 14306
rect 54574 14254 54626 14306
rect 15520 14086 15572 14138
rect 15624 14086 15676 14138
rect 15728 14086 15780 14138
rect 29827 14086 29879 14138
rect 29931 14086 29983 14138
rect 30035 14086 30087 14138
rect 44134 14086 44186 14138
rect 44238 14086 44290 14138
rect 44342 14086 44394 14138
rect 58441 14086 58493 14138
rect 58545 14086 58597 14138
rect 58649 14086 58701 14138
rect 5742 13918 5794 13970
rect 6638 13918 6690 13970
rect 6750 13918 6802 13970
rect 6862 13918 6914 13970
rect 9550 13918 9602 13970
rect 13806 13918 13858 13970
rect 15710 13918 15762 13970
rect 17390 13918 17442 13970
rect 18174 13918 18226 13970
rect 22542 13918 22594 13970
rect 23326 13918 23378 13970
rect 23774 13918 23826 13970
rect 25902 13918 25954 13970
rect 26798 13918 26850 13970
rect 27694 13918 27746 13970
rect 28478 13918 28530 13970
rect 29262 13918 29314 13970
rect 30718 13918 30770 13970
rect 34414 13918 34466 13970
rect 45054 13918 45106 13970
rect 49310 13918 49362 13970
rect 51214 13918 51266 13970
rect 55806 13918 55858 13970
rect 55918 13918 55970 13970
rect 2830 13806 2882 13858
rect 5966 13806 6018 13858
rect 12350 13806 12402 13858
rect 14702 13806 14754 13858
rect 15038 13806 15090 13858
rect 16718 13806 16770 13858
rect 21982 13806 22034 13858
rect 28702 13806 28754 13858
rect 28814 13806 28866 13858
rect 30046 13806 30098 13858
rect 36094 13806 36146 13858
rect 41582 13806 41634 13858
rect 44606 13806 44658 13858
rect 45502 13806 45554 13858
rect 48862 13806 48914 13858
rect 50318 13806 50370 13858
rect 51662 13806 51714 13858
rect 3950 13694 4002 13746
rect 4286 13694 4338 13746
rect 6190 13694 6242 13746
rect 7646 13694 7698 13746
rect 7870 13694 7922 13746
rect 8990 13694 9042 13746
rect 10446 13694 10498 13746
rect 11118 13694 11170 13746
rect 11342 13694 11394 13746
rect 11678 13694 11730 13746
rect 12686 13694 12738 13746
rect 16158 13694 16210 13746
rect 17614 13694 17666 13746
rect 18958 13694 19010 13746
rect 21198 13694 21250 13746
rect 25342 13694 25394 13746
rect 26686 13694 26738 13746
rect 26910 13694 26962 13746
rect 27806 13694 27858 13746
rect 27918 13694 27970 13746
rect 28366 13694 28418 13746
rect 30270 13694 30322 13746
rect 35758 13694 35810 13746
rect 36766 13694 36818 13746
rect 37438 13694 37490 13746
rect 40126 13694 40178 13746
rect 41358 13694 41410 13746
rect 42030 13694 42082 13746
rect 42254 13694 42306 13746
rect 44830 13694 44882 13746
rect 45726 13694 45778 13746
rect 48750 13694 48802 13746
rect 49870 13694 49922 13746
rect 52558 13694 52610 13746
rect 54350 13694 54402 13746
rect 54798 13694 54850 13746
rect 55358 13694 55410 13746
rect 56030 13694 56082 13746
rect 57598 13694 57650 13746
rect 1934 13582 1986 13634
rect 9662 13582 9714 13634
rect 10670 13582 10722 13634
rect 12798 13582 12850 13634
rect 18622 13582 18674 13634
rect 8766 13470 8818 13522
rect 10334 13470 10386 13522
rect 10782 13470 10834 13522
rect 18958 13582 19010 13634
rect 21086 13582 21138 13634
rect 24334 13582 24386 13634
rect 24670 13582 24722 13634
rect 25230 13582 25282 13634
rect 26462 13582 26514 13634
rect 29710 13582 29762 13634
rect 34750 13582 34802 13634
rect 34974 13582 35026 13634
rect 35870 13582 35922 13634
rect 37886 13582 37938 13634
rect 39566 13582 39618 13634
rect 42926 13582 42978 13634
rect 44158 13582 44210 13634
rect 44942 13582 44994 13634
rect 52894 13582 52946 13634
rect 57262 13582 57314 13634
rect 58158 13582 58210 13634
rect 15374 13470 15426 13522
rect 18734 13470 18786 13522
rect 21534 13470 21586 13522
rect 22206 13470 22258 13522
rect 26238 13470 26290 13522
rect 41022 13470 41074 13522
rect 45390 13470 45442 13522
rect 55022 13470 55074 13522
rect 8367 13302 8419 13354
rect 8471 13302 8523 13354
rect 8575 13302 8627 13354
rect 22674 13302 22726 13354
rect 22778 13302 22830 13354
rect 22882 13302 22934 13354
rect 36981 13302 37033 13354
rect 37085 13302 37137 13354
rect 37189 13302 37241 13354
rect 51288 13302 51340 13354
rect 51392 13302 51444 13354
rect 51496 13302 51548 13354
rect 2718 13134 2770 13186
rect 12238 13134 12290 13186
rect 17950 13134 18002 13186
rect 19630 13134 19682 13186
rect 28254 13134 28306 13186
rect 30942 13134 30994 13186
rect 46174 13134 46226 13186
rect 47294 13134 47346 13186
rect 48750 13134 48802 13186
rect 49086 13134 49138 13186
rect 49982 13134 50034 13186
rect 4398 13022 4450 13074
rect 4846 13022 4898 13074
rect 5966 13022 6018 13074
rect 8318 13022 8370 13074
rect 9886 13022 9938 13074
rect 10334 13022 10386 13074
rect 11118 13022 11170 13074
rect 14254 13022 14306 13074
rect 15374 13022 15426 13074
rect 16270 13022 16322 13074
rect 19294 13022 19346 13074
rect 20638 13022 20690 13074
rect 21422 13022 21474 13074
rect 22990 13022 23042 13074
rect 24782 13022 24834 13074
rect 28366 13022 28418 13074
rect 45166 13022 45218 13074
rect 46734 13022 46786 13074
rect 47630 13022 47682 13074
rect 50318 13022 50370 13074
rect 1934 12910 1986 12962
rect 4286 12910 4338 12962
rect 5070 12910 5122 12962
rect 8206 12910 8258 12962
rect 11006 12910 11058 12962
rect 11342 12910 11394 12962
rect 11678 12910 11730 12962
rect 12238 12910 12290 12962
rect 12574 12910 12626 12962
rect 14814 12910 14866 12962
rect 17614 12910 17666 12962
rect 18622 12910 18674 12962
rect 20190 12910 20242 12962
rect 21870 12910 21922 12962
rect 23326 12910 23378 12962
rect 26910 12910 26962 12962
rect 27246 12910 27298 12962
rect 28142 12910 28194 12962
rect 30606 12910 30658 12962
rect 31278 12910 31330 12962
rect 33294 12910 33346 12962
rect 35310 12910 35362 12962
rect 35870 12910 35922 12962
rect 37326 12910 37378 12962
rect 37550 12910 37602 12962
rect 37774 12910 37826 12962
rect 38558 12910 38610 12962
rect 39902 12910 39954 12962
rect 40350 12910 40402 12962
rect 45502 12910 45554 12962
rect 48078 12910 48130 12962
rect 48526 12910 48578 12962
rect 48974 12910 49026 12962
rect 9438 12798 9490 12850
rect 10670 12798 10722 12850
rect 15486 12798 15538 12850
rect 15934 12798 15986 12850
rect 16382 12798 16434 12850
rect 17054 12798 17106 12850
rect 17390 12798 17442 12850
rect 18510 12798 18562 12850
rect 22318 12798 22370 12850
rect 31390 12798 31442 12850
rect 33854 12798 33906 12850
rect 35758 12798 35810 12850
rect 37662 12798 37714 12850
rect 41246 12798 41298 12850
rect 3390 12686 3442 12738
rect 6302 12686 6354 12738
rect 6750 12686 6802 12738
rect 7198 12686 7250 12738
rect 13582 12686 13634 12738
rect 15262 12686 15314 12738
rect 16158 12686 16210 12738
rect 26462 12686 26514 12738
rect 29262 12686 29314 12738
rect 30830 12686 30882 12738
rect 34974 12686 35026 12738
rect 35534 12686 35586 12738
rect 41358 12686 41410 12738
rect 45838 12686 45890 12738
rect 46062 12686 46114 12738
rect 47518 12686 47570 12738
rect 48638 12686 48690 12738
rect 53118 13134 53170 13186
rect 55806 13134 55858 13186
rect 58046 13134 58098 13186
rect 51438 13022 51490 13074
rect 52894 13022 52946 13074
rect 54910 13022 54962 13074
rect 55470 13022 55522 13074
rect 56590 13022 56642 13074
rect 51102 12910 51154 12962
rect 51326 12910 51378 12962
rect 52670 12910 52722 12962
rect 53678 12910 53730 12962
rect 54462 12910 54514 12962
rect 55246 12910 55298 12962
rect 56030 12910 56082 12962
rect 56478 12910 56530 12962
rect 56702 12910 56754 12962
rect 57262 12910 57314 12962
rect 51550 12798 51602 12850
rect 51998 12798 52050 12850
rect 53342 12798 53394 12850
rect 57934 12798 57986 12850
rect 49870 12686 49922 12738
rect 50766 12686 50818 12738
rect 53230 12686 53282 12738
rect 54014 12686 54066 12738
rect 57038 12686 57090 12738
rect 57150 12686 57202 12738
rect 57486 12686 57538 12738
rect 58046 12686 58098 12738
rect 15520 12518 15572 12570
rect 15624 12518 15676 12570
rect 15728 12518 15780 12570
rect 29827 12518 29879 12570
rect 29931 12518 29983 12570
rect 30035 12518 30087 12570
rect 44134 12518 44186 12570
rect 44238 12518 44290 12570
rect 44342 12518 44394 12570
rect 58441 12518 58493 12570
rect 58545 12518 58597 12570
rect 58649 12518 58701 12570
rect 1934 12350 1986 12402
rect 9662 12350 9714 12402
rect 10558 12350 10610 12402
rect 11006 12350 11058 12402
rect 11454 12350 11506 12402
rect 12798 12350 12850 12402
rect 14142 12350 14194 12402
rect 15822 12350 15874 12402
rect 16382 12350 16434 12402
rect 18510 12350 18562 12402
rect 18734 12350 18786 12402
rect 18846 12350 18898 12402
rect 19630 12350 19682 12402
rect 22094 12350 22146 12402
rect 22542 12350 22594 12402
rect 22990 12350 23042 12402
rect 24670 12350 24722 12402
rect 29150 12350 29202 12402
rect 31278 12350 31330 12402
rect 36766 12350 36818 12402
rect 44382 12350 44434 12402
rect 45614 12350 45666 12402
rect 47518 12350 47570 12402
rect 47854 12350 47906 12402
rect 48078 12350 48130 12402
rect 50094 12350 50146 12402
rect 50766 12350 50818 12402
rect 52558 12350 52610 12402
rect 53006 12350 53058 12402
rect 55358 12350 55410 12402
rect 55582 12350 55634 12402
rect 55806 12350 55858 12402
rect 57598 12350 57650 12402
rect 2830 12238 2882 12290
rect 3838 12238 3890 12290
rect 5630 12238 5682 12290
rect 6190 12238 6242 12290
rect 15038 12238 15090 12290
rect 18398 12238 18450 12290
rect 19070 12238 19122 12290
rect 31054 12238 31106 12290
rect 35086 12238 35138 12290
rect 37438 12238 37490 12290
rect 47742 12238 47794 12290
rect 49646 12238 49698 12290
rect 51326 12238 51378 12290
rect 51662 12238 51714 12290
rect 52110 12238 52162 12290
rect 55694 12238 55746 12290
rect 57710 12238 57762 12290
rect 1598 12126 1650 12178
rect 1822 12126 1874 12178
rect 2494 12126 2546 12178
rect 3950 12126 4002 12178
rect 6974 12126 7026 12178
rect 12238 12126 12290 12178
rect 12574 12126 12626 12178
rect 14926 12126 14978 12178
rect 19182 12126 19234 12178
rect 23326 12126 23378 12178
rect 23550 12126 23602 12178
rect 25566 12126 25618 12178
rect 26126 12126 26178 12178
rect 28142 12126 28194 12178
rect 28366 12126 28418 12178
rect 29486 12126 29538 12178
rect 34190 12126 34242 12178
rect 35870 12126 35922 12178
rect 37998 12126 38050 12178
rect 41806 12126 41858 12178
rect 45166 12126 45218 12178
rect 48862 12126 48914 12178
rect 49422 12126 49474 12178
rect 51102 12126 51154 12178
rect 54238 12126 54290 12178
rect 54686 12126 54738 12178
rect 54798 12126 54850 12178
rect 54910 12126 54962 12178
rect 56702 12126 56754 12178
rect 57150 12126 57202 12178
rect 57374 12126 57426 12178
rect 57934 12126 57986 12178
rect 58158 12126 58210 12178
rect 8094 12014 8146 12066
rect 8542 12014 8594 12066
rect 8990 12014 9042 12066
rect 10110 12014 10162 12066
rect 12014 12014 12066 12066
rect 13694 12014 13746 12066
rect 17614 12014 17666 12066
rect 18062 12014 18114 12066
rect 21646 12014 21698 12066
rect 24110 12014 24162 12066
rect 27358 12014 27410 12066
rect 27918 12014 27970 12066
rect 31166 12014 31218 12066
rect 42030 12014 42082 12066
rect 43038 12014 43090 12066
rect 44718 12014 44770 12066
rect 46958 12014 47010 12066
rect 49310 12014 49362 12066
rect 51550 12014 51602 12066
rect 53790 12014 53842 12066
rect 57262 12014 57314 12066
rect 7310 11902 7362 11954
rect 14478 11902 14530 11954
rect 44942 11902 44994 11954
rect 49086 11902 49138 11954
rect 8367 11734 8419 11786
rect 8471 11734 8523 11786
rect 8575 11734 8627 11786
rect 22674 11734 22726 11786
rect 22778 11734 22830 11786
rect 22882 11734 22934 11786
rect 36981 11734 37033 11786
rect 37085 11734 37137 11786
rect 37189 11734 37241 11786
rect 51288 11734 51340 11786
rect 51392 11734 51444 11786
rect 51496 11734 51548 11786
rect 2270 11566 2322 11618
rect 2718 11566 2770 11618
rect 6974 11566 7026 11618
rect 9662 11566 9714 11618
rect 11790 11566 11842 11618
rect 21870 11566 21922 11618
rect 22094 11566 22146 11618
rect 30158 11566 30210 11618
rect 4510 11454 4562 11506
rect 4958 11454 5010 11506
rect 5742 11454 5794 11506
rect 10782 11454 10834 11506
rect 11230 11454 11282 11506
rect 12574 11454 12626 11506
rect 13022 11454 13074 11506
rect 13694 11454 13746 11506
rect 14142 11454 14194 11506
rect 14590 11454 14642 11506
rect 18958 11454 19010 11506
rect 26238 11454 26290 11506
rect 26798 11454 26850 11506
rect 31166 11454 31218 11506
rect 39454 11454 39506 11506
rect 40014 11454 40066 11506
rect 41918 11454 41970 11506
rect 44942 11454 44994 11506
rect 45950 11454 46002 11506
rect 47518 11454 47570 11506
rect 48302 11454 48354 11506
rect 49086 11454 49138 11506
rect 50318 11454 50370 11506
rect 50654 11454 50706 11506
rect 51774 11454 51826 11506
rect 53566 11454 53618 11506
rect 54014 11454 54066 11506
rect 57486 11454 57538 11506
rect 2494 11342 2546 11394
rect 6862 11342 6914 11394
rect 7870 11342 7922 11394
rect 9438 11342 9490 11394
rect 11454 11342 11506 11394
rect 19294 11342 19346 11394
rect 20750 11342 20802 11394
rect 22318 11342 22370 11394
rect 23326 11342 23378 11394
rect 23774 11342 23826 11394
rect 23998 11342 24050 11394
rect 27134 11342 27186 11394
rect 30382 11342 30434 11394
rect 38670 11342 38722 11394
rect 39006 11342 39058 11394
rect 40238 11342 40290 11394
rect 41694 11342 41746 11394
rect 44718 11342 44770 11394
rect 45278 11342 45330 11394
rect 51662 11342 51714 11394
rect 55134 11342 55186 11394
rect 55918 11342 55970 11394
rect 56254 11342 56306 11394
rect 56702 11342 56754 11394
rect 2046 11230 2098 11282
rect 7086 11230 7138 11282
rect 9102 11230 9154 11282
rect 15262 11230 15314 11282
rect 19630 11230 19682 11282
rect 22542 11230 22594 11282
rect 22990 11230 23042 11282
rect 23102 11230 23154 11282
rect 25790 11230 25842 11282
rect 28142 11230 28194 11282
rect 30046 11230 30098 11282
rect 31278 11230 31330 11282
rect 32958 11230 33010 11282
rect 33182 11230 33234 11282
rect 39902 11230 39954 11282
rect 44270 11230 44322 11282
rect 45166 11230 45218 11282
rect 46846 11230 46898 11282
rect 46958 11230 47010 11282
rect 52110 11230 52162 11282
rect 54910 11230 54962 11282
rect 57822 11230 57874 11282
rect 3166 11118 3218 11170
rect 3502 11118 3554 11170
rect 3950 11118 4002 11170
rect 6190 11118 6242 11170
rect 9998 11118 10050 11170
rect 11678 11118 11730 11170
rect 15710 11118 15762 11170
rect 19518 11118 19570 11170
rect 21422 11118 21474 11170
rect 28478 11118 28530 11170
rect 29822 11118 29874 11170
rect 38222 11118 38274 11170
rect 40686 11118 40738 11170
rect 42926 11118 42978 11170
rect 46286 11118 46338 11170
rect 47182 11118 47234 11170
rect 48638 11118 48690 11170
rect 49534 11118 49586 11170
rect 54686 11118 54738 11170
rect 55470 11118 55522 11170
rect 56366 11118 56418 11170
rect 57374 11118 57426 11170
rect 57598 11118 57650 11170
rect 15520 10950 15572 11002
rect 15624 10950 15676 11002
rect 15728 10950 15780 11002
rect 29827 10950 29879 11002
rect 29931 10950 29983 11002
rect 30035 10950 30087 11002
rect 44134 10950 44186 11002
rect 44238 10950 44290 11002
rect 44342 10950 44394 11002
rect 58441 10950 58493 11002
rect 58545 10950 58597 11002
rect 58649 10950 58701 11002
rect 2270 10782 2322 10834
rect 15486 10782 15538 10834
rect 24110 10782 24162 10834
rect 24670 10782 24722 10834
rect 25902 10782 25954 10834
rect 26574 10782 26626 10834
rect 27358 10782 27410 10834
rect 29150 10782 29202 10834
rect 29934 10782 29986 10834
rect 30494 10782 30546 10834
rect 38334 10782 38386 10834
rect 55246 10782 55298 10834
rect 55806 10782 55858 10834
rect 56030 10782 56082 10834
rect 56142 10782 56194 10834
rect 3054 10670 3106 10722
rect 9662 10670 9714 10722
rect 12126 10670 12178 10722
rect 12574 10670 12626 10722
rect 13470 10670 13522 10722
rect 13582 10670 13634 10722
rect 14142 10670 14194 10722
rect 16606 10670 16658 10722
rect 17390 10670 17442 10722
rect 19294 10670 19346 10722
rect 21646 10670 21698 10722
rect 21870 10670 21922 10722
rect 29486 10670 29538 10722
rect 32286 10670 32338 10722
rect 34974 10670 35026 10722
rect 36318 10670 36370 10722
rect 39342 10670 39394 10722
rect 40014 10670 40066 10722
rect 41246 10670 41298 10722
rect 42030 10670 42082 10722
rect 46398 10670 46450 10722
rect 46622 10670 46674 10722
rect 47294 10670 47346 10722
rect 48862 10670 48914 10722
rect 49758 10670 49810 10722
rect 49982 10670 50034 10722
rect 51774 10670 51826 10722
rect 55582 10670 55634 10722
rect 2942 10558 2994 10610
rect 5630 10558 5682 10610
rect 7198 10558 7250 10610
rect 7422 10558 7474 10610
rect 10670 10558 10722 10610
rect 11230 10558 11282 10610
rect 13022 10558 13074 10610
rect 14366 10558 14418 10610
rect 14590 10558 14642 10610
rect 14702 10558 14754 10610
rect 15374 10558 15426 10610
rect 15710 10558 15762 10610
rect 16270 10558 16322 10610
rect 17614 10558 17666 10610
rect 20750 10558 20802 10610
rect 21086 10558 21138 10610
rect 22430 10558 22482 10610
rect 22878 10558 22930 10610
rect 23326 10558 23378 10610
rect 25454 10558 25506 10610
rect 26350 10558 26402 10610
rect 26574 10558 26626 10610
rect 26910 10558 26962 10610
rect 28142 10558 28194 10610
rect 28366 10558 28418 10610
rect 31502 10558 31554 10610
rect 31726 10558 31778 10610
rect 34862 10558 34914 10610
rect 39118 10558 39170 10610
rect 39566 10558 39618 10610
rect 40126 10558 40178 10610
rect 41582 10558 41634 10610
rect 41918 10558 41970 10610
rect 42254 10558 42306 10610
rect 43038 10558 43090 10610
rect 43486 10558 43538 10610
rect 45054 10558 45106 10610
rect 47406 10558 47458 10610
rect 47854 10558 47906 10610
rect 49310 10558 49362 10610
rect 51998 10558 52050 10610
rect 52894 10558 52946 10610
rect 56926 10558 56978 10610
rect 3054 10446 3106 10498
rect 4958 10446 5010 10498
rect 5854 10446 5906 10498
rect 13806 10446 13858 10498
rect 14478 10446 14530 10498
rect 28814 10446 28866 10498
rect 39790 10446 39842 10498
rect 40910 10446 40962 10498
rect 45278 10446 45330 10498
rect 46734 10446 46786 10498
rect 47630 10446 47682 10498
rect 49534 10446 49586 10498
rect 50430 10446 50482 10498
rect 54686 10446 54738 10498
rect 2830 10334 2882 10386
rect 8318 10334 8370 10386
rect 9886 10334 9938 10386
rect 10222 10334 10274 10386
rect 10782 10334 10834 10386
rect 12798 10334 12850 10386
rect 16046 10334 16098 10386
rect 16718 10334 16770 10386
rect 16830 10334 16882 10386
rect 17838 10334 17890 10386
rect 18062 10334 18114 10386
rect 18510 10334 18562 10386
rect 21982 10334 22034 10386
rect 23438 10334 23490 10386
rect 29374 10334 29426 10386
rect 37662 10334 37714 10386
rect 38782 10334 38834 10386
rect 48078 10334 48130 10386
rect 54238 10334 54290 10386
rect 54686 10334 54738 10386
rect 55134 10334 55186 10386
rect 57934 10334 57986 10386
rect 8367 10166 8419 10218
rect 8471 10166 8523 10218
rect 8575 10166 8627 10218
rect 22674 10166 22726 10218
rect 22778 10166 22830 10218
rect 22882 10166 22934 10218
rect 36981 10166 37033 10218
rect 37085 10166 37137 10218
rect 37189 10166 37241 10218
rect 51288 10166 51340 10218
rect 51392 10166 51444 10218
rect 51496 10166 51548 10218
rect 4622 9998 4674 10050
rect 6638 9998 6690 10050
rect 9438 9998 9490 10050
rect 13918 9998 13970 10050
rect 19966 9998 20018 10050
rect 27022 9998 27074 10050
rect 28030 9998 28082 10050
rect 47966 9998 48018 10050
rect 49646 9998 49698 10050
rect 4510 9886 4562 9938
rect 6750 9886 6802 9938
rect 11566 9886 11618 9938
rect 13694 9886 13746 9938
rect 14254 9886 14306 9938
rect 15374 9886 15426 9938
rect 18286 9886 18338 9938
rect 27582 9886 27634 9938
rect 28030 9886 28082 9938
rect 30718 9886 30770 9938
rect 38446 9886 38498 9938
rect 41806 9886 41858 9938
rect 42926 9886 42978 9938
rect 46958 9886 47010 9938
rect 49982 9886 50034 9938
rect 1934 9774 1986 9826
rect 3950 9774 4002 9826
rect 4174 9774 4226 9826
rect 6078 9774 6130 9826
rect 6302 9774 6354 9826
rect 7646 9774 7698 9826
rect 9102 9774 9154 9826
rect 9998 9774 10050 9826
rect 10446 9774 10498 9826
rect 15710 9774 15762 9826
rect 16158 9774 16210 9826
rect 18958 9774 19010 9826
rect 22654 9774 22706 9826
rect 24670 9774 24722 9826
rect 30270 9774 30322 9826
rect 31278 9774 31330 9826
rect 31614 9774 31666 9826
rect 34302 9774 34354 9826
rect 35198 9774 35250 9826
rect 38110 9774 38162 9826
rect 40126 9774 40178 9826
rect 40462 9774 40514 9826
rect 42590 9774 42642 9826
rect 45054 9774 45106 9826
rect 46734 9774 46786 9826
rect 48190 9774 48242 9826
rect 48414 9774 48466 9826
rect 48526 9774 48578 9826
rect 49086 9774 49138 9826
rect 49310 9774 49362 9826
rect 56030 9774 56082 9826
rect 56478 9774 56530 9826
rect 2494 9662 2546 9714
rect 7758 9662 7810 9714
rect 8878 9662 8930 9714
rect 11230 9662 11282 9714
rect 17838 9662 17890 9714
rect 18846 9662 18898 9714
rect 23214 9662 23266 9714
rect 26350 9662 26402 9714
rect 32846 9662 32898 9714
rect 34190 9662 34242 9714
rect 36430 9662 36482 9714
rect 38334 9662 38386 9714
rect 39342 9662 39394 9714
rect 40350 9662 40402 9714
rect 42366 9662 42418 9714
rect 46510 9662 46562 9714
rect 49534 9662 49586 9714
rect 54910 9662 54962 9714
rect 58158 9662 58210 9714
rect 8094 9550 8146 9602
rect 12574 9550 12626 9602
rect 14702 9550 14754 9602
rect 24110 9550 24162 9602
rect 27022 9550 27074 9602
rect 30606 9550 30658 9602
rect 30830 9550 30882 9602
rect 42814 9550 42866 9602
rect 42926 9550 42978 9602
rect 43486 9550 43538 9602
rect 48078 9550 48130 9602
rect 54574 9550 54626 9602
rect 15520 9382 15572 9434
rect 15624 9382 15676 9434
rect 15728 9382 15780 9434
rect 29827 9382 29879 9434
rect 29931 9382 29983 9434
rect 30035 9382 30087 9434
rect 44134 9382 44186 9434
rect 44238 9382 44290 9434
rect 44342 9382 44394 9434
rect 58441 9382 58493 9434
rect 58545 9382 58597 9434
rect 58649 9382 58701 9434
rect 5070 9214 5122 9266
rect 7534 9214 7586 9266
rect 7982 9214 8034 9266
rect 9662 9214 9714 9266
rect 10110 9214 10162 9266
rect 21646 9214 21698 9266
rect 39454 9214 39506 9266
rect 41022 9214 41074 9266
rect 47070 9214 47122 9266
rect 50430 9214 50482 9266
rect 3726 9102 3778 9154
rect 3838 9102 3890 9154
rect 4510 9102 4562 9154
rect 4846 9102 4898 9154
rect 5182 9102 5234 9154
rect 7086 9102 7138 9154
rect 10670 9102 10722 9154
rect 11230 9102 11282 9154
rect 13806 9102 13858 9154
rect 14702 9102 14754 9154
rect 15598 9102 15650 9154
rect 17726 9102 17778 9154
rect 18062 9102 18114 9154
rect 19182 9102 19234 9154
rect 22542 9102 22594 9154
rect 24446 9102 24498 9154
rect 25790 9102 25842 9154
rect 26686 9102 26738 9154
rect 27358 9102 27410 9154
rect 37102 9102 37154 9154
rect 37214 9102 37266 9154
rect 41582 9102 41634 9154
rect 42590 9102 42642 9154
rect 43598 9102 43650 9154
rect 44606 9102 44658 9154
rect 46398 9102 46450 9154
rect 48750 9102 48802 9154
rect 48974 9102 49026 9154
rect 57374 9102 57426 9154
rect 2718 8990 2770 9042
rect 3390 8990 3442 9042
rect 4062 8990 4114 9042
rect 4398 8990 4450 9042
rect 9998 8990 10050 9042
rect 10334 8990 10386 9042
rect 10782 8990 10834 9042
rect 14478 8990 14530 9042
rect 18286 8990 18338 9042
rect 18510 8990 18562 9042
rect 18734 8990 18786 9042
rect 19070 8990 19122 9042
rect 21982 8990 22034 9042
rect 23662 8990 23714 9042
rect 25230 8990 25282 9042
rect 25454 8990 25506 9042
rect 26014 8990 26066 9042
rect 26462 8990 26514 9042
rect 27582 8990 27634 9042
rect 28030 8990 28082 9042
rect 41134 8990 41186 9042
rect 41918 8990 41970 9042
rect 43038 8990 43090 9042
rect 44718 8990 44770 9042
rect 47630 8990 47682 9042
rect 48078 8990 48130 9042
rect 48190 8990 48242 9042
rect 50766 8990 50818 9042
rect 50990 8990 51042 9042
rect 52894 8990 52946 9042
rect 53230 8990 53282 9042
rect 55358 8990 55410 9042
rect 56478 8990 56530 9042
rect 57598 8990 57650 9042
rect 2046 8878 2098 8930
rect 3950 8878 4002 8930
rect 5742 8878 5794 8930
rect 8542 8878 8594 8930
rect 8990 8878 9042 8930
rect 13358 8878 13410 8930
rect 15150 8878 15202 8930
rect 18622 8878 18674 8930
rect 26574 8878 26626 8930
rect 31054 8878 31106 8930
rect 51326 8878 51378 8930
rect 52110 8878 52162 8930
rect 53566 8878 53618 8930
rect 55246 8878 55298 8930
rect 57710 8878 57762 8930
rect 4510 8766 4562 8818
rect 6526 8766 6578 8818
rect 6862 8766 6914 8818
rect 7646 8766 7698 8818
rect 8990 8766 9042 8818
rect 10670 8766 10722 8818
rect 28366 8766 28418 8818
rect 37214 8766 37266 8818
rect 47518 8766 47570 8818
rect 47854 8766 47906 8818
rect 49086 8766 49138 8818
rect 8367 8598 8419 8650
rect 8471 8598 8523 8650
rect 8575 8598 8627 8650
rect 22674 8598 22726 8650
rect 22778 8598 22830 8650
rect 22882 8598 22934 8650
rect 36981 8598 37033 8650
rect 37085 8598 37137 8650
rect 37189 8598 37241 8650
rect 51288 8598 51340 8650
rect 51392 8598 51444 8650
rect 51496 8598 51548 8650
rect 10782 8430 10834 8482
rect 25902 8430 25954 8482
rect 35086 8430 35138 8482
rect 37214 8430 37266 8482
rect 39230 8430 39282 8482
rect 43150 8430 43202 8482
rect 47854 8430 47906 8482
rect 48302 8430 48354 8482
rect 2046 8318 2098 8370
rect 3950 8318 4002 8370
rect 4846 8318 4898 8370
rect 5742 8318 5794 8370
rect 10334 8318 10386 8370
rect 11230 8318 11282 8370
rect 12910 8318 12962 8370
rect 14926 8318 14978 8370
rect 20190 8318 20242 8370
rect 21310 8318 21362 8370
rect 24558 8318 24610 8370
rect 31838 8318 31890 8370
rect 33518 8318 33570 8370
rect 37438 8318 37490 8370
rect 37774 8318 37826 8370
rect 42142 8318 42194 8370
rect 45950 8318 46002 8370
rect 49086 8318 49138 8370
rect 50318 8318 50370 8370
rect 50654 8318 50706 8370
rect 56478 8318 56530 8370
rect 57150 8318 57202 8370
rect 3166 8206 3218 8258
rect 6414 8206 6466 8258
rect 7422 8206 7474 8258
rect 7982 8206 8034 8258
rect 8206 8206 8258 8258
rect 9438 8206 9490 8258
rect 9774 8206 9826 8258
rect 10446 8206 10498 8258
rect 11342 8206 11394 8258
rect 12462 8206 12514 8258
rect 13470 8206 13522 8258
rect 13918 8206 13970 8258
rect 19854 8206 19906 8258
rect 21534 8206 21586 8258
rect 21870 8206 21922 8258
rect 22318 8206 22370 8258
rect 22878 8206 22930 8258
rect 25006 8206 25058 8258
rect 26014 8206 26066 8258
rect 26462 8206 26514 8258
rect 26910 8206 26962 8258
rect 27134 8206 27186 8258
rect 27806 8206 27858 8258
rect 28030 8206 28082 8258
rect 29710 8206 29762 8258
rect 31054 8206 31106 8258
rect 32734 8206 32786 8258
rect 33406 8206 33458 8258
rect 34078 8206 34130 8258
rect 35870 8206 35922 8258
rect 37998 8206 38050 8258
rect 39342 8206 39394 8258
rect 40686 8206 40738 8258
rect 41806 8206 41858 8258
rect 42478 8206 42530 8258
rect 42702 8206 42754 8258
rect 43486 8206 43538 8258
rect 45054 8206 45106 8258
rect 46398 8206 46450 8258
rect 47630 8206 47682 8258
rect 48078 8206 48130 8258
rect 48414 8206 48466 8258
rect 48750 8206 48802 8258
rect 50878 8206 50930 8258
rect 53790 8206 53842 8258
rect 54798 8206 54850 8258
rect 57262 8206 57314 8258
rect 57710 8206 57762 8258
rect 2382 8094 2434 8146
rect 6302 8094 6354 8146
rect 6750 8094 6802 8146
rect 7310 8094 7362 8146
rect 8878 8094 8930 8146
rect 9214 8094 9266 8146
rect 14142 8094 14194 8146
rect 15486 8094 15538 8146
rect 15598 8094 15650 8146
rect 15710 8094 15762 8146
rect 20526 8094 20578 8146
rect 23886 8094 23938 8146
rect 25454 8094 25506 8146
rect 27358 8094 27410 8146
rect 27470 8094 27522 8146
rect 28142 8094 28194 8146
rect 28590 8094 28642 8146
rect 29150 8094 29202 8146
rect 29374 8094 29426 8146
rect 31166 8094 31218 8146
rect 31614 8094 31666 8146
rect 32510 8094 32562 8146
rect 33630 8094 33682 8146
rect 34974 8094 35026 8146
rect 35534 8094 35586 8146
rect 37438 8094 37490 8146
rect 42254 8094 42306 8146
rect 43374 8094 43426 8146
rect 44046 8094 44098 8146
rect 44830 8094 44882 8146
rect 45166 8094 45218 8146
rect 46846 8094 46898 8146
rect 51550 8094 51602 8146
rect 54014 8094 54066 8146
rect 54686 8094 54738 8146
rect 2494 7982 2546 8034
rect 2718 7982 2770 8034
rect 6078 7982 6130 8034
rect 7646 7982 7698 8034
rect 7758 7982 7810 8034
rect 13694 7982 13746 8034
rect 13806 7982 13858 8034
rect 15262 7982 15314 8034
rect 15374 7982 15426 8034
rect 25902 7982 25954 8034
rect 29598 7982 29650 8034
rect 31390 7982 31442 8034
rect 32174 7982 32226 8034
rect 33070 7982 33122 8034
rect 35086 7982 35138 8034
rect 35646 7982 35698 8034
rect 45838 7982 45890 8034
rect 46062 7982 46114 8034
rect 46734 7982 46786 8034
rect 48974 7982 49026 8034
rect 52894 7982 52946 8034
rect 15520 7814 15572 7866
rect 15624 7814 15676 7866
rect 15728 7814 15780 7866
rect 29827 7814 29879 7866
rect 29931 7814 29983 7866
rect 30035 7814 30087 7866
rect 44134 7814 44186 7866
rect 44238 7814 44290 7866
rect 44342 7814 44394 7866
rect 58441 7814 58493 7866
rect 58545 7814 58597 7866
rect 58649 7814 58701 7866
rect 1822 7646 1874 7698
rect 5294 7646 5346 7698
rect 5630 7646 5682 7698
rect 7534 7646 7586 7698
rect 7982 7646 8034 7698
rect 8430 7646 8482 7698
rect 9438 7646 9490 7698
rect 9662 7646 9714 7698
rect 18174 7646 18226 7698
rect 24670 7646 24722 7698
rect 34862 7646 34914 7698
rect 41022 7646 41074 7698
rect 43598 7646 43650 7698
rect 45278 7646 45330 7698
rect 46062 7646 46114 7698
rect 46398 7646 46450 7698
rect 47182 7646 47234 7698
rect 48862 7646 48914 7698
rect 3390 7534 3442 7586
rect 3838 7534 3890 7586
rect 12126 7534 12178 7586
rect 14030 7534 14082 7586
rect 25678 7534 25730 7586
rect 25790 7534 25842 7586
rect 27470 7534 27522 7586
rect 30830 7534 30882 7586
rect 34190 7534 34242 7586
rect 38782 7534 38834 7586
rect 40910 7534 40962 7586
rect 41246 7534 41298 7586
rect 42142 7534 42194 7586
rect 44718 7534 44770 7586
rect 45054 7534 45106 7586
rect 45838 7534 45890 7586
rect 46958 7534 47010 7586
rect 2830 7422 2882 7474
rect 4062 7422 4114 7474
rect 4398 7422 4450 7474
rect 6190 7422 6242 7474
rect 7086 7422 7138 7474
rect 9774 7422 9826 7474
rect 10334 7422 10386 7474
rect 10558 7422 10610 7474
rect 11230 7422 11282 7474
rect 11902 7422 11954 7474
rect 12574 7422 12626 7474
rect 12910 7422 12962 7474
rect 14590 7422 14642 7474
rect 15374 7422 15426 7474
rect 17838 7422 17890 7474
rect 18174 7422 18226 7474
rect 18510 7422 18562 7474
rect 20190 7422 20242 7474
rect 20414 7422 20466 7474
rect 21086 7422 21138 7474
rect 26014 7422 26066 7474
rect 27694 7422 27746 7474
rect 28254 7422 28306 7474
rect 28926 7422 28978 7474
rect 29934 7422 29986 7474
rect 30270 7422 30322 7474
rect 34526 7422 34578 7474
rect 34750 7422 34802 7474
rect 40126 7422 40178 7474
rect 42030 7422 42082 7474
rect 43710 7422 43762 7474
rect 45726 7422 45778 7474
rect 46286 7422 46338 7474
rect 46622 7422 46674 7474
rect 46846 7422 46898 7474
rect 57150 7422 57202 7474
rect 58046 7422 58098 7474
rect 2382 7310 2434 7362
rect 6526 7310 6578 7362
rect 12238 7310 12290 7362
rect 13358 7310 13410 7362
rect 15934 7310 15986 7362
rect 45390 7310 45442 7362
rect 48078 7310 48130 7362
rect 56814 7310 56866 7362
rect 57598 7310 57650 7362
rect 7198 7198 7250 7250
rect 7758 7198 7810 7250
rect 25230 7198 25282 7250
rect 29038 7198 29090 7250
rect 33966 7198 34018 7250
rect 39118 7198 39170 7250
rect 57934 7198 57986 7250
rect 8367 7030 8419 7082
rect 8471 7030 8523 7082
rect 8575 7030 8627 7082
rect 22674 7030 22726 7082
rect 22778 7030 22830 7082
rect 22882 7030 22934 7082
rect 36981 7030 37033 7082
rect 37085 7030 37137 7082
rect 37189 7030 37241 7082
rect 51288 7030 51340 7082
rect 51392 7030 51444 7082
rect 51496 7030 51548 7082
rect 3278 6862 3330 6914
rect 3614 6862 3666 6914
rect 4398 6862 4450 6914
rect 4846 6862 4898 6914
rect 16158 6862 16210 6914
rect 27582 6862 27634 6914
rect 27918 6862 27970 6914
rect 35646 6862 35698 6914
rect 43150 6862 43202 6914
rect 43934 6862 43986 6914
rect 44270 6862 44322 6914
rect 46846 6862 46898 6914
rect 52782 6862 52834 6914
rect 2718 6750 2770 6802
rect 4398 6750 4450 6802
rect 4734 6750 4786 6802
rect 6526 6750 6578 6802
rect 7758 6750 7810 6802
rect 9998 6750 10050 6802
rect 15598 6750 15650 6802
rect 17502 6750 17554 6802
rect 24222 6750 24274 6802
rect 28142 6750 28194 6802
rect 35422 6750 35474 6802
rect 42702 6750 42754 6802
rect 51102 6750 51154 6802
rect 55022 6750 55074 6802
rect 1710 6638 1762 6690
rect 3838 6638 3890 6690
rect 5742 6638 5794 6690
rect 6414 6638 6466 6690
rect 7534 6638 7586 6690
rect 15934 6638 15986 6690
rect 16382 6638 16434 6690
rect 17390 6638 17442 6690
rect 18174 6638 18226 6690
rect 18510 6638 18562 6690
rect 24110 6638 24162 6690
rect 33070 6638 33122 6690
rect 33966 6638 34018 6690
rect 34638 6638 34690 6690
rect 35198 6638 35250 6690
rect 38222 6638 38274 6690
rect 39230 6638 39282 6690
rect 40910 6638 40962 6690
rect 41246 6638 41298 6690
rect 42030 6638 42082 6690
rect 42814 6638 42866 6690
rect 44270 6638 44322 6690
rect 44830 6638 44882 6690
rect 46062 6638 46114 6690
rect 46734 6638 46786 6690
rect 47182 6638 47234 6690
rect 48526 6638 48578 6690
rect 48750 6638 48802 6690
rect 48974 6638 49026 6690
rect 50766 6638 50818 6690
rect 54910 6638 54962 6690
rect 55358 6638 55410 6690
rect 57038 6638 57090 6690
rect 57374 6638 57426 6690
rect 6190 6526 6242 6578
rect 18062 6526 18114 6578
rect 25006 6526 25058 6578
rect 25118 6526 25170 6578
rect 32734 6526 32786 6578
rect 33630 6526 33682 6578
rect 33742 6526 33794 6578
rect 39006 6526 39058 6578
rect 52670 6526 52722 6578
rect 7870 6414 7922 6466
rect 23886 6414 23938 6466
rect 24782 6414 24834 6466
rect 32398 6414 32450 6466
rect 32846 6414 32898 6466
rect 50094 6414 50146 6466
rect 51998 6414 52050 6466
rect 52782 6414 52834 6466
rect 15520 6246 15572 6298
rect 15624 6246 15676 6298
rect 15728 6246 15780 6298
rect 29827 6246 29879 6298
rect 29931 6246 29983 6298
rect 30035 6246 30087 6298
rect 44134 6246 44186 6298
rect 44238 6246 44290 6298
rect 44342 6246 44394 6298
rect 58441 6246 58493 6298
rect 58545 6246 58597 6298
rect 58649 6246 58701 6298
rect 1822 6078 1874 6130
rect 3502 6078 3554 6130
rect 4734 6078 4786 6130
rect 5070 6078 5122 6130
rect 5518 6078 5570 6130
rect 6638 6078 6690 6130
rect 6974 6078 7026 6130
rect 7758 6078 7810 6130
rect 8430 6078 8482 6130
rect 19294 6078 19346 6130
rect 21758 6078 21810 6130
rect 25342 6078 25394 6130
rect 28254 6078 28306 6130
rect 28814 6078 28866 6130
rect 36990 6078 37042 6130
rect 37550 6078 37602 6130
rect 38222 6078 38274 6130
rect 39902 6078 39954 6130
rect 40126 6078 40178 6130
rect 42142 6078 42194 6130
rect 50654 6078 50706 6130
rect 51326 6078 51378 6130
rect 51662 6078 51714 6130
rect 52222 6078 52274 6130
rect 54014 6078 54066 6130
rect 56142 6078 56194 6130
rect 18398 5966 18450 6018
rect 19070 5966 19122 6018
rect 21422 5966 21474 6018
rect 27358 5966 27410 6018
rect 33294 5966 33346 6018
rect 38446 5966 38498 6018
rect 43038 5966 43090 6018
rect 48078 5966 48130 6018
rect 50094 5966 50146 6018
rect 50990 5966 51042 6018
rect 51102 5966 51154 6018
rect 52110 5966 52162 6018
rect 2606 5854 2658 5906
rect 8206 5854 8258 5906
rect 8318 5854 8370 5906
rect 8766 5854 8818 5906
rect 10222 5854 10274 5906
rect 10446 5854 10498 5906
rect 10670 5854 10722 5906
rect 18846 5854 18898 5906
rect 19406 5854 19458 5906
rect 21646 5854 21698 5906
rect 22094 5854 22146 5906
rect 22430 5854 22482 5906
rect 27022 5854 27074 5906
rect 27806 5854 27858 5906
rect 31726 5854 31778 5906
rect 31950 5854 32002 5906
rect 32398 5854 32450 5906
rect 34974 5854 35026 5906
rect 35198 5854 35250 5906
rect 35646 5854 35698 5906
rect 37886 5854 37938 5906
rect 38334 5854 38386 5906
rect 39790 5854 39842 5906
rect 42030 5854 42082 5906
rect 42814 5854 42866 5906
rect 46846 5854 46898 5906
rect 47070 5854 47122 5906
rect 47630 5854 47682 5906
rect 48862 5854 48914 5906
rect 48974 5854 49026 5906
rect 49086 5854 49138 5906
rect 49198 5854 49250 5906
rect 49534 5854 49586 5906
rect 50318 5854 50370 5906
rect 54014 5854 54066 5906
rect 54350 5854 54402 5906
rect 55694 5854 55746 5906
rect 56926 5854 56978 5906
rect 58046 5854 58098 5906
rect 2382 5742 2434 5794
rect 3838 5742 3890 5794
rect 6078 5742 6130 5794
rect 10558 5742 10610 5794
rect 35086 5742 35138 5794
rect 42702 5742 42754 5794
rect 53902 5742 53954 5794
rect 55246 5742 55298 5794
rect 55470 5742 55522 5794
rect 2942 5630 2994 5682
rect 5070 5630 5122 5682
rect 6078 5630 6130 5682
rect 18510 5630 18562 5682
rect 27022 5630 27074 5682
rect 32174 5630 32226 5682
rect 32510 5630 32562 5682
rect 33070 5630 33122 5682
rect 33406 5630 33458 5682
rect 52222 5630 52274 5682
rect 8367 5462 8419 5514
rect 8471 5462 8523 5514
rect 8575 5462 8627 5514
rect 22674 5462 22726 5514
rect 22778 5462 22830 5514
rect 22882 5462 22934 5514
rect 36981 5462 37033 5514
rect 37085 5462 37137 5514
rect 37189 5462 37241 5514
rect 51288 5462 51340 5514
rect 51392 5462 51444 5514
rect 51496 5462 51548 5514
rect 4734 5294 4786 5346
rect 11678 5294 11730 5346
rect 18958 5294 19010 5346
rect 28254 5294 28306 5346
rect 28478 5294 28530 5346
rect 29598 5294 29650 5346
rect 35086 5294 35138 5346
rect 35758 5294 35810 5346
rect 38334 5294 38386 5346
rect 47070 5294 47122 5346
rect 49198 5294 49250 5346
rect 2270 5182 2322 5234
rect 2718 5182 2770 5234
rect 3166 5182 3218 5234
rect 7310 5182 7362 5234
rect 8206 5182 8258 5234
rect 10782 5182 10834 5234
rect 12686 5182 12738 5234
rect 13806 5182 13858 5234
rect 19294 5182 19346 5234
rect 22542 5182 22594 5234
rect 23998 5182 24050 5234
rect 27246 5182 27298 5234
rect 30606 5182 30658 5234
rect 31502 5182 31554 5234
rect 34414 5182 34466 5234
rect 34526 5182 34578 5234
rect 34862 5182 34914 5234
rect 35870 5182 35922 5234
rect 37662 5182 37714 5234
rect 38558 5182 38610 5234
rect 41582 5182 41634 5234
rect 43374 5182 43426 5234
rect 48750 5182 48802 5234
rect 49422 5182 49474 5234
rect 49758 5182 49810 5234
rect 50878 5182 50930 5234
rect 51326 5182 51378 5234
rect 55470 5182 55522 5234
rect 1822 5070 1874 5122
rect 3726 5070 3778 5122
rect 4174 5070 4226 5122
rect 4846 5070 4898 5122
rect 5742 5070 5794 5122
rect 6190 5070 6242 5122
rect 8094 5070 8146 5122
rect 8318 5070 8370 5122
rect 8766 5070 8818 5122
rect 9214 5070 9266 5122
rect 10894 5070 10946 5122
rect 13582 5070 13634 5122
rect 15598 5070 15650 5122
rect 16382 5070 16434 5122
rect 20190 5070 20242 5122
rect 20526 5070 20578 5122
rect 20638 5070 20690 5122
rect 23326 5070 23378 5122
rect 23662 5070 23714 5122
rect 25790 5070 25842 5122
rect 27806 5070 27858 5122
rect 28142 5070 28194 5122
rect 29710 5070 29762 5122
rect 30830 5070 30882 5122
rect 39454 5070 39506 5122
rect 39790 5070 39842 5122
rect 40686 5070 40738 5122
rect 43598 5070 43650 5122
rect 43822 5070 43874 5122
rect 45278 5070 45330 5122
rect 45614 5070 45666 5122
rect 46734 5070 46786 5122
rect 48302 5070 48354 5122
rect 54574 5070 54626 5122
rect 55582 5070 55634 5122
rect 57486 5070 57538 5122
rect 57710 5070 57762 5122
rect 4958 4958 5010 5010
rect 9550 4958 9602 5010
rect 13918 4958 13970 5010
rect 15822 4958 15874 5010
rect 19182 4958 19234 5010
rect 25566 4958 25618 5010
rect 29150 4958 29202 5010
rect 29374 4958 29426 5010
rect 39902 4958 39954 5010
rect 12798 4846 12850 4898
rect 16718 4846 16770 4898
rect 20750 4846 20802 4898
rect 27134 4846 27186 4898
rect 27358 4846 27410 4898
rect 28142 4846 28194 4898
rect 29262 4846 29314 4898
rect 35422 4846 35474 4898
rect 37998 4846 38050 4898
rect 39118 4846 39170 4898
rect 40014 4846 40066 4898
rect 44942 4846 44994 4898
rect 49646 4846 49698 4898
rect 49870 4846 49922 4898
rect 50430 4846 50482 4898
rect 15520 4678 15572 4730
rect 15624 4678 15676 4730
rect 15728 4678 15780 4730
rect 29827 4678 29879 4730
rect 29931 4678 29983 4730
rect 30035 4678 30087 4730
rect 44134 4678 44186 4730
rect 44238 4678 44290 4730
rect 44342 4678 44394 4730
rect 58441 4678 58493 4730
rect 58545 4678 58597 4730
rect 58649 4678 58701 4730
rect 2046 4510 2098 4562
rect 2494 4510 2546 4562
rect 3166 4510 3218 4562
rect 4398 4510 4450 4562
rect 4958 4510 5010 4562
rect 5182 4510 5234 4562
rect 5294 4510 5346 4562
rect 5630 4510 5682 4562
rect 6638 4510 6690 4562
rect 9550 4510 9602 4562
rect 9774 4510 9826 4562
rect 13470 4510 13522 4562
rect 19966 4510 20018 4562
rect 23998 4510 24050 4562
rect 24334 4510 24386 4562
rect 25230 4510 25282 4562
rect 25454 4510 25506 4562
rect 27694 4510 27746 4562
rect 28478 4510 28530 4562
rect 36318 4510 36370 4562
rect 40350 4510 40402 4562
rect 44494 4510 44546 4562
rect 47966 4510 48018 4562
rect 48974 4510 49026 4562
rect 55806 4510 55858 4562
rect 56030 4510 56082 4562
rect 58046 4510 58098 4562
rect 8206 4398 8258 4450
rect 9886 4398 9938 4450
rect 12910 4398 12962 4450
rect 14478 4398 14530 4450
rect 16158 4398 16210 4450
rect 16382 4398 16434 4450
rect 18062 4398 18114 4450
rect 19518 4398 19570 4450
rect 19742 4398 19794 4450
rect 20078 4398 20130 4450
rect 20638 4398 20690 4450
rect 21422 4398 21474 4450
rect 22766 4398 22818 4450
rect 24110 4398 24162 4450
rect 25566 4398 25618 4450
rect 26686 4398 26738 4450
rect 30606 4398 30658 4450
rect 32510 4398 32562 4450
rect 33294 4398 33346 4450
rect 37326 4398 37378 4450
rect 38670 4398 38722 4450
rect 41358 4398 41410 4450
rect 45166 4398 45218 4450
rect 47406 4398 47458 4450
rect 47742 4398 47794 4450
rect 51550 4398 51602 4450
rect 1822 4286 1874 4338
rect 4622 4286 4674 4338
rect 6078 4286 6130 4338
rect 6302 4286 6354 4338
rect 7534 4286 7586 4338
rect 7982 4286 8034 4338
rect 10558 4286 10610 4338
rect 11006 4286 11058 4338
rect 12014 4286 12066 4338
rect 12462 4286 12514 4338
rect 13246 4286 13298 4338
rect 13358 4286 13410 4338
rect 13806 4286 13858 4338
rect 17950 4286 18002 4338
rect 18734 4286 18786 4338
rect 20974 4286 21026 4338
rect 22430 4286 22482 4338
rect 22878 4286 22930 4338
rect 23774 4286 23826 4338
rect 24670 4286 24722 4338
rect 25902 4286 25954 4338
rect 27134 4286 27186 4338
rect 28366 4286 28418 4338
rect 28590 4286 28642 4338
rect 29038 4286 29090 4338
rect 30830 4286 30882 4338
rect 31950 4286 32002 4338
rect 32286 4286 32338 4338
rect 33070 4286 33122 4338
rect 37438 4286 37490 4338
rect 39230 4286 39282 4338
rect 41246 4286 41298 4338
rect 41582 4286 41634 4338
rect 42590 4286 42642 4338
rect 43822 4286 43874 4338
rect 44158 4286 44210 4338
rect 49310 4286 49362 4338
rect 49534 4286 49586 4338
rect 51102 4286 51154 4338
rect 55470 4286 55522 4338
rect 57598 4286 57650 4338
rect 57822 4286 57874 4338
rect 3614 4174 3666 4226
rect 4062 4174 4114 4226
rect 11454 4174 11506 4226
rect 14254 4174 14306 4226
rect 26014 4174 26066 4226
rect 26798 4174 26850 4226
rect 31166 4174 31218 4226
rect 33182 4174 33234 4226
rect 39006 4174 39058 4226
rect 48078 4174 48130 4226
rect 50206 4174 50258 4226
rect 50654 4174 50706 4226
rect 55918 4174 55970 4226
rect 3390 4062 3442 4114
rect 3614 4062 3666 4114
rect 4062 4062 4114 4114
rect 19070 4062 19122 4114
rect 20974 4062 21026 4114
rect 21870 4062 21922 4114
rect 23438 4062 23490 4114
rect 23774 4062 23826 4114
rect 26462 4062 26514 4114
rect 27358 4062 27410 4114
rect 36654 4062 36706 4114
rect 8367 3894 8419 3946
rect 8471 3894 8523 3946
rect 8575 3894 8627 3946
rect 22674 3894 22726 3946
rect 22778 3894 22830 3946
rect 22882 3894 22934 3946
rect 36981 3894 37033 3946
rect 37085 3894 37137 3946
rect 37189 3894 37241 3946
rect 51288 3894 51340 3946
rect 51392 3894 51444 3946
rect 51496 3894 51548 3946
rect 6862 3726 6914 3778
rect 13470 3726 13522 3778
rect 21870 3726 21922 3778
rect 22206 3726 22258 3778
rect 32958 3726 33010 3778
rect 36542 3726 36594 3778
rect 36878 3726 36930 3778
rect 56814 3726 56866 3778
rect 57038 3726 57090 3778
rect 2830 3614 2882 3666
rect 3502 3614 3554 3666
rect 3950 3614 4002 3666
rect 4734 3614 4786 3666
rect 7198 3614 7250 3666
rect 13246 3614 13298 3666
rect 23662 3614 23714 3666
rect 25678 3614 25730 3666
rect 32286 3614 32338 3666
rect 32846 3614 32898 3666
rect 41246 3614 41298 3666
rect 42030 3614 42082 3666
rect 43934 3614 43986 3666
rect 44718 3614 44770 3666
rect 46846 3614 46898 3666
rect 47630 3614 47682 3666
rect 48190 3614 48242 3666
rect 56590 3614 56642 3666
rect 57486 3614 57538 3666
rect 1710 3502 1762 3554
rect 6302 3502 6354 3554
rect 6526 3502 6578 3554
rect 13134 3502 13186 3554
rect 21646 3502 21698 3554
rect 24558 3502 24610 3554
rect 24894 3502 24946 3554
rect 25118 3502 25170 3554
rect 25566 3502 25618 3554
rect 32622 3502 32674 3554
rect 37550 3502 37602 3554
rect 41470 3502 41522 3554
rect 42366 3502 42418 3554
rect 44830 3502 44882 3554
rect 48526 3502 48578 3554
rect 55582 3502 55634 3554
rect 57934 3502 57986 3554
rect 4286 3390 4338 3442
rect 6750 3390 6802 3442
rect 23774 3390 23826 3442
rect 24670 3390 24722 3442
rect 25790 3390 25842 3442
rect 37662 3390 37714 3442
rect 41918 3390 41970 3442
rect 42702 3390 42754 3442
rect 48974 3390 49026 3442
rect 56254 3390 56306 3442
rect 57598 3390 57650 3442
rect 57822 3390 57874 3442
rect 15520 3110 15572 3162
rect 15624 3110 15676 3162
rect 15728 3110 15780 3162
rect 29827 3110 29879 3162
rect 29931 3110 29983 3162
rect 30035 3110 30087 3162
rect 44134 3110 44186 3162
rect 44238 3110 44290 3162
rect 44342 3110 44394 3162
rect 58441 3110 58493 3162
rect 58545 3110 58597 3162
rect 58649 3110 58701 3162
<< metal2 >>
rect 9856 29200 9968 30000
rect 29792 29200 29904 30000
rect 49728 29200 49840 30000
rect 5516 28308 5572 28318
rect 2156 26516 2212 26526
rect 1484 26404 1540 26414
rect 1260 26068 1316 26078
rect 1260 13188 1316 26012
rect 1260 13122 1316 13132
rect 1484 13076 1540 26348
rect 2156 26290 2212 26460
rect 2156 26238 2158 26290
rect 2210 26238 2212 26290
rect 1708 25506 1764 25518
rect 1708 25454 1710 25506
rect 1762 25454 1764 25506
rect 1708 24724 1764 25454
rect 1708 24658 1764 24668
rect 1708 24498 1764 24510
rect 1708 24446 1710 24498
rect 1762 24446 1764 24498
rect 1708 23266 1764 24446
rect 2156 23492 2212 26238
rect 5516 26290 5572 28252
rect 7980 26516 8036 26526
rect 7980 26402 8036 26460
rect 7980 26350 7982 26402
rect 8034 26350 8036 26402
rect 7980 26338 8036 26350
rect 8204 26402 8260 26414
rect 8204 26350 8206 26402
rect 8258 26350 8260 26402
rect 5516 26238 5518 26290
rect 5570 26238 5572 26290
rect 5068 26178 5124 26190
rect 5068 26126 5070 26178
rect 5122 26126 5124 26178
rect 4060 26066 4116 26078
rect 4060 26014 4062 26066
rect 4114 26014 4116 26066
rect 4060 25732 4116 26014
rect 4060 25666 4116 25676
rect 3052 25618 3108 25630
rect 3052 25566 3054 25618
rect 3106 25566 3108 25618
rect 3052 25396 3108 25566
rect 2492 24724 2548 24734
rect 2492 24722 2660 24724
rect 2492 24670 2494 24722
rect 2546 24670 2660 24722
rect 2492 24668 2660 24670
rect 2492 24658 2548 24668
rect 2156 23426 2212 23436
rect 2268 23714 2324 23726
rect 2268 23662 2270 23714
rect 2322 23662 2324 23714
rect 1708 23214 1710 23266
rect 1762 23214 1764 23266
rect 1708 21812 1764 23214
rect 2268 23156 2324 23662
rect 2268 23090 2324 23100
rect 2492 23154 2548 23166
rect 2492 23102 2494 23154
rect 2546 23102 2548 23154
rect 1820 22930 1876 22942
rect 1820 22878 1822 22930
rect 1874 22878 1876 22930
rect 1820 22820 1876 22878
rect 1820 22754 1876 22764
rect 1708 21746 1764 21756
rect 2380 22372 2436 22382
rect 2492 22372 2548 23102
rect 2604 22932 2660 24668
rect 3052 23938 3108 25340
rect 4844 25284 4900 25294
rect 3052 23886 3054 23938
rect 3106 23886 3108 23938
rect 2940 23268 2996 23278
rect 2940 23174 2996 23212
rect 2604 22866 2660 22876
rect 2716 23042 2772 23054
rect 2716 22990 2718 23042
rect 2770 22990 2772 23042
rect 2380 22370 2548 22372
rect 2380 22318 2382 22370
rect 2434 22318 2548 22370
rect 2380 22316 2548 22318
rect 2716 22820 2772 22990
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21140 1764 21534
rect 1708 21074 1764 21084
rect 1820 20804 1876 20814
rect 2380 20804 2436 22316
rect 2716 22258 2772 22764
rect 2716 22206 2718 22258
rect 2770 22206 2772 22258
rect 2716 22194 2772 22206
rect 1820 20802 2436 20804
rect 1820 20750 1822 20802
rect 1874 20750 2436 20802
rect 1820 20748 2436 20750
rect 2604 21812 2660 21822
rect 2604 20802 2660 21756
rect 2604 20750 2606 20802
rect 2658 20750 2660 20802
rect 1708 19348 1764 19358
rect 1708 19234 1764 19292
rect 1708 19182 1710 19234
rect 1762 19182 1764 19234
rect 1708 19170 1764 19182
rect 1820 18116 1876 20748
rect 2604 20738 2660 20750
rect 2716 21474 2772 21486
rect 2716 21422 2718 21474
rect 2770 21422 2772 21474
rect 2268 20578 2324 20590
rect 2268 20526 2270 20578
rect 2322 20526 2324 20578
rect 2268 20356 2324 20526
rect 2268 20290 2324 20300
rect 2716 20244 2772 21422
rect 2940 20690 2996 20702
rect 2940 20638 2942 20690
rect 2994 20638 2996 20690
rect 2940 20356 2996 20638
rect 2940 20290 2996 20300
rect 2716 20178 2772 20188
rect 2156 20130 2212 20142
rect 2156 20078 2158 20130
rect 2210 20078 2212 20130
rect 2044 20020 2100 20030
rect 2044 19926 2100 19964
rect 2156 20020 2212 20078
rect 2940 20020 2996 20030
rect 2156 20018 2996 20020
rect 2156 19966 2942 20018
rect 2994 19966 2996 20018
rect 2156 19964 2996 19966
rect 2044 19796 2100 19806
rect 1932 19794 2100 19796
rect 1932 19742 2046 19794
rect 2098 19742 2100 19794
rect 1932 19740 2100 19742
rect 1932 18340 1988 19740
rect 2044 19730 2100 19740
rect 2156 18674 2212 19964
rect 2940 19954 2996 19964
rect 2492 19796 2548 19806
rect 2156 18622 2158 18674
rect 2210 18622 2212 18674
rect 2156 18610 2212 18622
rect 2268 19122 2324 19134
rect 2268 19070 2270 19122
rect 2322 19070 2324 19122
rect 1932 18274 1988 18284
rect 2044 18450 2100 18462
rect 2044 18398 2046 18450
rect 2098 18398 2100 18450
rect 1820 18060 1988 18116
rect 1820 17666 1876 17678
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 17556 1876 17614
rect 1708 15876 1764 15886
rect 1484 13010 1540 13020
rect 1596 15874 1764 15876
rect 1596 15822 1710 15874
rect 1762 15822 1764 15874
rect 1596 15820 1764 15822
rect 1596 15764 1652 15820
rect 1708 15810 1764 15820
rect 1596 12178 1652 15708
rect 1820 14868 1876 17500
rect 1932 15316 1988 18060
rect 2044 17780 2100 18398
rect 2268 17892 2324 19070
rect 2044 17714 2100 17724
rect 2156 17836 2324 17892
rect 2492 18338 2548 19740
rect 2828 18452 2884 18462
rect 2828 18358 2884 18396
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2044 16772 2100 16782
rect 2044 16678 2100 16716
rect 1932 15250 1988 15260
rect 1820 14802 1876 14812
rect 2044 15202 2100 15214
rect 2044 15150 2046 15202
rect 2098 15150 2100 15202
rect 1820 14644 1876 14654
rect 1596 12126 1598 12178
rect 1650 12126 1652 12178
rect 1596 12114 1652 12126
rect 1708 14306 1764 14318
rect 1708 14254 1710 14306
rect 1762 14254 1764 14306
rect 1708 13972 1764 14254
rect 1708 7476 1764 13916
rect 1820 12404 1876 14588
rect 2044 13972 2100 15150
rect 2156 14868 2212 17836
rect 2268 17666 2324 17678
rect 2268 17614 2270 17666
rect 2322 17614 2324 17666
rect 2268 17108 2324 17614
rect 2268 17042 2324 17052
rect 2268 16884 2324 16894
rect 2492 16884 2548 18286
rect 2940 17780 2996 17790
rect 2940 17686 2996 17724
rect 3052 17556 3108 23886
rect 3164 24722 3220 24734
rect 3164 24670 3166 24722
rect 3218 24670 3220 24722
rect 3164 23380 3220 24670
rect 3724 24722 3780 24734
rect 3724 24670 3726 24722
rect 3778 24670 3780 24722
rect 3276 24052 3332 24062
rect 3276 23958 3332 23996
rect 3164 23324 3668 23380
rect 3612 23042 3668 23324
rect 3724 23268 3780 24670
rect 4732 24724 4788 24734
rect 4620 23828 4676 23838
rect 4620 23734 4676 23772
rect 3724 23154 3780 23212
rect 4732 23268 4788 24668
rect 4732 23202 4788 23212
rect 3724 23102 3726 23154
rect 3778 23102 3780 23154
rect 3724 23090 3780 23102
rect 3836 23156 3892 23166
rect 4620 23156 4676 23166
rect 3892 23100 4004 23156
rect 3836 23090 3892 23100
rect 3612 22990 3614 23042
rect 3666 22990 3668 23042
rect 3388 22148 3444 22158
rect 3612 22148 3668 22990
rect 3388 22146 3668 22148
rect 3388 22094 3390 22146
rect 3442 22094 3668 22146
rect 3388 22092 3668 22094
rect 3388 22082 3444 22092
rect 3388 21812 3444 21822
rect 3164 21756 3388 21812
rect 3164 20188 3220 21756
rect 3388 21718 3444 21756
rect 3500 21588 3556 21598
rect 3836 21588 3892 21598
rect 3500 21494 3556 21532
rect 3612 21586 3892 21588
rect 3612 21534 3838 21586
rect 3890 21534 3892 21586
rect 3612 21532 3892 21534
rect 3388 21364 3444 21374
rect 3612 21364 3668 21532
rect 3836 21522 3892 21532
rect 3388 21362 3668 21364
rect 3388 21310 3390 21362
rect 3442 21310 3668 21362
rect 3388 21308 3668 21310
rect 3388 21298 3444 21308
rect 3948 20804 4004 23100
rect 3724 20748 4004 20804
rect 4060 22932 4116 22942
rect 3276 20692 3332 20702
rect 3276 20598 3332 20636
rect 3612 20356 3668 20366
rect 3164 20132 3444 20188
rect 3164 20020 3220 20030
rect 3164 19926 3220 19964
rect 2324 16828 2548 16884
rect 2716 17500 3108 17556
rect 2268 16658 2324 16828
rect 2268 16606 2270 16658
rect 2322 16606 2324 16658
rect 2268 16436 2324 16606
rect 2268 16370 2324 16380
rect 2492 16658 2548 16670
rect 2492 16606 2494 16658
rect 2546 16606 2548 16658
rect 2492 16324 2548 16606
rect 2716 16658 2772 17500
rect 3276 17444 3332 20132
rect 3388 20020 3444 20132
rect 3388 19954 3444 19964
rect 3500 19236 3556 19246
rect 2940 17388 3332 17444
rect 3388 17554 3444 17566
rect 3388 17502 3390 17554
rect 3442 17502 3444 17554
rect 2940 16772 2996 17388
rect 3388 17220 3444 17502
rect 3388 17154 3444 17164
rect 3052 17108 3108 17118
rect 3108 17052 3332 17108
rect 3052 17042 3108 17052
rect 2940 16706 2996 16716
rect 3164 16660 3220 16670
rect 2716 16606 2718 16658
rect 2770 16606 2772 16658
rect 2716 16548 2772 16606
rect 2716 16482 2772 16492
rect 3052 16658 3220 16660
rect 3052 16606 3166 16658
rect 3218 16606 3220 16658
rect 3052 16604 3220 16606
rect 2492 16258 2548 16268
rect 2268 16098 2324 16110
rect 3052 16100 3108 16604
rect 3164 16594 3220 16604
rect 2268 16046 2270 16098
rect 2322 16046 2324 16098
rect 2268 15428 2324 16046
rect 2268 15362 2324 15372
rect 2380 16098 3108 16100
rect 2380 16046 3054 16098
rect 3106 16046 3108 16098
rect 2380 16044 3108 16046
rect 2380 15314 2436 16044
rect 3052 16034 3108 16044
rect 3164 16436 3220 16446
rect 2604 15428 2660 15438
rect 2604 15334 2660 15372
rect 2828 15428 2884 15438
rect 2380 15262 2382 15314
rect 2434 15262 2436 15314
rect 2380 15250 2436 15262
rect 2716 15316 2772 15326
rect 2156 14802 2212 14812
rect 2604 15092 2660 15102
rect 2604 14530 2660 15036
rect 2604 14478 2606 14530
rect 2658 14478 2660 14530
rect 2604 14466 2660 14478
rect 2268 14418 2324 14430
rect 2268 14366 2270 14418
rect 2322 14366 2324 14418
rect 2268 14084 2324 14366
rect 2716 14308 2772 15260
rect 2828 15148 2884 15372
rect 3052 15316 3108 15326
rect 3164 15316 3220 16380
rect 3052 15314 3220 15316
rect 3052 15262 3054 15314
rect 3106 15262 3220 15314
rect 3052 15260 3220 15262
rect 3052 15250 3108 15260
rect 2828 15092 3108 15148
rect 2940 14532 2996 14542
rect 2940 14438 2996 14476
rect 2716 14306 2884 14308
rect 2716 14254 2718 14306
rect 2770 14254 2884 14306
rect 2716 14252 2884 14254
rect 2716 14242 2772 14252
rect 2268 14018 2324 14028
rect 2044 13916 2212 13972
rect 2156 13860 2212 13916
rect 2716 13860 2772 13870
rect 2156 13804 2324 13860
rect 1932 13636 1988 13646
rect 1932 13542 1988 13580
rect 1932 12962 1988 12974
rect 1932 12910 1934 12962
rect 1986 12910 1988 12962
rect 1932 12852 1988 12910
rect 1932 12786 1988 12796
rect 2156 12852 2212 12862
rect 1932 12404 1988 12414
rect 1820 12402 1988 12404
rect 1820 12350 1934 12402
rect 1986 12350 1988 12402
rect 1820 12348 1988 12350
rect 1932 12338 1988 12348
rect 1820 12178 1876 12190
rect 1820 12126 1822 12178
rect 1874 12126 1876 12178
rect 1820 7698 1876 12126
rect 2156 12180 2212 12796
rect 2044 11396 2100 11406
rect 2044 11282 2100 11340
rect 2044 11230 2046 11282
rect 2098 11230 2100 11282
rect 1932 10276 1988 10286
rect 1932 9826 1988 10220
rect 1932 9774 1934 9826
rect 1986 9774 1988 9826
rect 1932 9716 1988 9774
rect 1932 9650 1988 9660
rect 2044 8930 2100 11230
rect 2044 8878 2046 8930
rect 2098 8878 2100 8930
rect 2044 8866 2100 8878
rect 2044 8372 2100 8382
rect 2156 8372 2212 12124
rect 2268 11956 2324 13804
rect 2268 11890 2324 11900
rect 2380 13636 2436 13646
rect 2268 11620 2324 11630
rect 2380 11620 2436 13580
rect 2716 13188 2772 13804
rect 2828 13860 2884 14252
rect 2828 13858 2996 13860
rect 2828 13806 2830 13858
rect 2882 13806 2996 13858
rect 2828 13804 2996 13806
rect 2828 13794 2884 13804
rect 2940 13412 2996 13804
rect 3052 13524 3108 15092
rect 3052 13458 3108 13468
rect 3164 14868 3220 14878
rect 2716 13186 2884 13188
rect 2716 13134 2718 13186
rect 2770 13134 2884 13186
rect 2716 13132 2884 13134
rect 2716 13122 2772 13132
rect 2828 12292 2884 13132
rect 2716 12290 2884 12292
rect 2716 12238 2830 12290
rect 2882 12238 2884 12290
rect 2716 12236 2884 12238
rect 2268 11618 2380 11620
rect 2268 11566 2270 11618
rect 2322 11566 2380 11618
rect 2268 11564 2380 11566
rect 2268 11554 2324 11564
rect 2380 11526 2436 11564
rect 2492 12178 2548 12190
rect 2492 12126 2494 12178
rect 2546 12126 2548 12178
rect 2492 11732 2548 12126
rect 2492 11394 2548 11676
rect 2716 11618 2772 12236
rect 2828 12226 2884 12236
rect 2828 12068 2884 12078
rect 2940 12068 2996 13356
rect 3164 12516 3220 14812
rect 3164 12450 3220 12460
rect 2884 12012 2996 12068
rect 2828 12002 2884 12012
rect 2940 11844 2996 11854
rect 2716 11566 2718 11618
rect 2770 11566 2772 11618
rect 2716 11554 2772 11566
rect 2828 11788 2940 11844
rect 3276 11844 3332 17052
rect 3500 16996 3556 19180
rect 3612 19234 3668 20300
rect 3612 19182 3614 19234
rect 3666 19182 3668 19234
rect 3612 19170 3668 19182
rect 3388 16940 3556 16996
rect 3612 18564 3668 18574
rect 3724 18564 3780 20748
rect 3948 19908 4004 19918
rect 3948 19234 4004 19852
rect 3948 19182 3950 19234
rect 4002 19182 4004 19234
rect 3948 19170 4004 19182
rect 3612 18562 3780 18564
rect 3612 18510 3614 18562
rect 3666 18510 3780 18562
rect 3612 18508 3780 18510
rect 3948 18564 4004 18574
rect 3612 17780 3668 18508
rect 3948 18470 4004 18508
rect 3836 18452 3892 18462
rect 3836 18358 3892 18396
rect 3612 17554 3668 17724
rect 3612 17502 3614 17554
rect 3666 17502 3668 17554
rect 3388 16322 3444 16940
rect 3388 16270 3390 16322
rect 3442 16270 3444 16322
rect 3388 16212 3444 16270
rect 3388 16146 3444 16156
rect 3500 16772 3556 16782
rect 3500 15428 3556 16716
rect 3500 15362 3556 15372
rect 3612 15148 3668 17502
rect 3724 17778 3780 17790
rect 3724 17726 3726 17778
rect 3778 17726 3780 17778
rect 3724 16884 3780 17726
rect 3724 16818 3780 16828
rect 3612 15092 3780 15148
rect 3612 14196 3668 14206
rect 3500 13524 3556 13534
rect 3388 12738 3444 12750
rect 3388 12686 3390 12738
rect 3442 12686 3444 12738
rect 3388 12180 3444 12686
rect 3388 12114 3444 12124
rect 3276 11788 3444 11844
rect 2492 11342 2494 11394
rect 2546 11342 2548 11394
rect 2268 10836 2324 10846
rect 2268 10742 2324 10780
rect 2492 9714 2548 11342
rect 2828 10386 2884 11788
rect 2940 11778 2996 11788
rect 3052 11396 3108 11406
rect 3052 10722 3108 11340
rect 3052 10670 3054 10722
rect 3106 10670 3108 10722
rect 3052 10658 3108 10670
rect 3164 11170 3220 11182
rect 3164 11118 3166 11170
rect 3218 11118 3220 11170
rect 2940 10612 2996 10622
rect 2940 10518 2996 10556
rect 2828 10334 2830 10386
rect 2882 10334 2884 10386
rect 2828 10322 2884 10334
rect 3052 10498 3108 10510
rect 3052 10446 3054 10498
rect 3106 10446 3108 10498
rect 3052 9828 3108 10446
rect 2492 9662 2494 9714
rect 2546 9662 2548 9714
rect 2492 8708 2548 9662
rect 2492 8642 2548 8652
rect 2604 9716 2660 9726
rect 2044 8370 2212 8372
rect 2044 8318 2046 8370
rect 2098 8318 2212 8370
rect 2044 8316 2212 8318
rect 2044 8306 2100 8316
rect 2380 8148 2436 8158
rect 1820 7646 1822 7698
rect 1874 7646 1876 7698
rect 1820 7634 1876 7646
rect 2268 8092 2380 8148
rect 1708 7420 1876 7476
rect 1708 6692 1764 6702
rect 1708 6598 1764 6636
rect 1820 6356 1876 7420
rect 2268 7140 2324 8092
rect 2380 8054 2436 8092
rect 2492 8034 2548 8046
rect 2492 7982 2494 8034
rect 2546 7982 2548 8034
rect 2492 7812 2548 7982
rect 2380 7364 2436 7374
rect 2492 7364 2548 7756
rect 2380 7362 2548 7364
rect 2380 7310 2382 7362
rect 2434 7310 2548 7362
rect 2380 7308 2548 7310
rect 2380 7298 2436 7308
rect 2604 7252 2660 9660
rect 2716 9042 2772 9054
rect 2716 8990 2718 9042
rect 2770 8990 2772 9042
rect 2716 8596 2772 8990
rect 2772 8540 2884 8596
rect 2716 8530 2772 8540
rect 2716 8036 2772 8046
rect 2716 7942 2772 7980
rect 2828 7700 2884 8540
rect 3052 7924 3108 9772
rect 3164 8260 3220 11118
rect 3388 9268 3444 11788
rect 3500 11396 3556 13468
rect 3612 11508 3668 14140
rect 3724 13748 3780 15092
rect 3948 14530 4004 14542
rect 3948 14478 3950 14530
rect 4002 14478 4004 14530
rect 3948 14420 4004 14478
rect 3948 14354 4004 14364
rect 3948 13748 4004 13758
rect 3724 13746 4004 13748
rect 3724 13694 3950 13746
rect 4002 13694 4004 13746
rect 3724 13692 4004 13694
rect 3836 13412 3892 13422
rect 3836 12290 3892 13356
rect 3836 12238 3838 12290
rect 3890 12238 3892 12290
rect 3836 12226 3892 12238
rect 3948 12740 4004 13692
rect 3948 12180 4004 12684
rect 3948 11508 4004 12124
rect 3612 11452 3780 11508
rect 3500 11340 3668 11396
rect 3500 11172 3556 11182
rect 3500 11078 3556 11116
rect 3612 10052 3668 11340
rect 3388 9202 3444 9212
rect 3500 9996 3668 10052
rect 3388 9042 3444 9054
rect 3388 8990 3390 9042
rect 3442 8990 3444 9042
rect 3388 8932 3444 8990
rect 3500 9044 3556 9996
rect 3500 8978 3556 8988
rect 3612 9380 3668 9390
rect 3388 8866 3444 8876
rect 3612 8820 3668 9324
rect 3724 9154 3780 11452
rect 3948 11170 4004 11452
rect 3948 11118 3950 11170
rect 4002 11118 4004 11170
rect 3948 10948 4004 11118
rect 3948 10882 4004 10892
rect 4060 10836 4116 22876
rect 4396 22370 4452 22382
rect 4396 22318 4398 22370
rect 4450 22318 4452 22370
rect 4284 19348 4340 19358
rect 4172 18450 4228 18462
rect 4172 18398 4174 18450
rect 4226 18398 4228 18450
rect 4172 16882 4228 18398
rect 4284 17778 4340 19292
rect 4396 18674 4452 22318
rect 4620 22258 4676 23100
rect 4844 22930 4900 25228
rect 4844 22878 4846 22930
rect 4898 22878 4900 22930
rect 4844 22866 4900 22878
rect 4956 24722 5012 24734
rect 4956 24670 4958 24722
rect 5010 24670 5012 24722
rect 4956 22932 5012 24670
rect 5068 23714 5124 26126
rect 5068 23662 5070 23714
rect 5122 23662 5124 23714
rect 5068 23044 5124 23662
rect 5068 22978 5124 22988
rect 5180 25282 5236 25294
rect 5180 25230 5182 25282
rect 5234 25230 5236 25282
rect 5180 23828 5236 25230
rect 4956 22866 5012 22876
rect 5180 22820 5236 23772
rect 5404 24722 5460 24734
rect 5404 24670 5406 24722
rect 5458 24670 5460 24722
rect 5404 23156 5460 24670
rect 5404 23090 5460 23100
rect 4620 22206 4622 22258
rect 4674 22206 4676 22258
rect 4620 22194 4676 22206
rect 5068 22764 5236 22820
rect 5516 22820 5572 26238
rect 6860 26290 6916 26302
rect 6860 26238 6862 26290
rect 6914 26238 6916 26290
rect 5964 26180 6020 26190
rect 5964 26086 6020 26124
rect 5852 25732 5908 25742
rect 5852 25618 5908 25676
rect 5852 25566 5854 25618
rect 5906 25566 5908 25618
rect 5852 25554 5908 25566
rect 6860 25620 6916 26238
rect 7196 26290 7252 26302
rect 7196 26238 7198 26290
rect 7250 26238 7252 26290
rect 7196 25732 7252 26238
rect 7308 26292 7364 26302
rect 7308 26198 7364 26236
rect 7644 26290 7700 26302
rect 7644 26238 7646 26290
rect 7698 26238 7700 26290
rect 7196 25666 7252 25676
rect 7644 26068 7700 26238
rect 6860 25554 6916 25564
rect 7532 25620 7588 25630
rect 6972 25506 7028 25518
rect 6972 25454 6974 25506
rect 7026 25454 7028 25506
rect 6972 25396 7028 25454
rect 6972 25330 7028 25340
rect 7196 25506 7252 25518
rect 7196 25454 7198 25506
rect 7250 25454 7252 25506
rect 6300 25282 6356 25294
rect 6300 25230 6302 25282
rect 6354 25230 6356 25282
rect 5628 24836 5684 24846
rect 5628 24742 5684 24780
rect 5740 23826 5796 23838
rect 5740 23774 5742 23826
rect 5794 23774 5796 23826
rect 5740 23156 5796 23774
rect 5964 23156 6020 23166
rect 5740 23154 6020 23156
rect 5740 23102 5966 23154
rect 6018 23102 6020 23154
rect 5740 23100 6020 23102
rect 5628 22820 5684 22830
rect 5516 22764 5628 22820
rect 4956 21924 5012 21934
rect 4396 18622 4398 18674
rect 4450 18622 4452 18674
rect 4396 18452 4452 18622
rect 4396 18386 4452 18396
rect 4508 21588 4564 21598
rect 4508 20916 4564 21532
rect 4956 21026 5012 21868
rect 4956 20974 4958 21026
rect 5010 20974 5012 21026
rect 4956 20962 5012 20974
rect 4508 18450 4564 20860
rect 4620 20804 4676 20814
rect 4620 20690 4676 20748
rect 4620 20638 4622 20690
rect 4674 20638 4676 20690
rect 4620 20130 4676 20638
rect 4732 20802 4788 20814
rect 4732 20750 4734 20802
rect 4786 20750 4788 20802
rect 4732 20692 4788 20750
rect 4732 20626 4788 20636
rect 4620 20078 4622 20130
rect 4674 20078 4676 20130
rect 4620 20066 4676 20078
rect 4844 19908 4900 19918
rect 4844 19814 4900 19852
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 4284 17726 4286 17778
rect 4338 17726 4340 17778
rect 4284 17714 4340 17726
rect 4508 17444 4564 18398
rect 4508 17378 4564 17388
rect 4620 19124 4676 19134
rect 4620 16996 4676 19068
rect 5068 19012 5124 22764
rect 5628 22754 5684 22764
rect 5964 22260 6020 23100
rect 6300 23044 6356 25230
rect 6636 25282 6692 25294
rect 6636 25230 6638 25282
rect 6690 25230 6692 25282
rect 6412 24722 6468 24734
rect 6412 24670 6414 24722
rect 6466 24670 6468 24722
rect 6412 24052 6468 24670
rect 6636 24724 6692 25230
rect 7196 25060 7252 25454
rect 7532 25060 7588 25564
rect 7644 25284 7700 26012
rect 7644 25218 7700 25228
rect 7756 25506 7812 25518
rect 7756 25454 7758 25506
rect 7810 25454 7812 25506
rect 7532 25004 7700 25060
rect 7196 24994 7252 25004
rect 6636 24658 6692 24668
rect 7644 24722 7700 25004
rect 7644 24670 7646 24722
rect 7698 24670 7700 24722
rect 7196 24610 7252 24622
rect 7196 24558 7198 24610
rect 7250 24558 7252 24610
rect 6636 24500 6692 24510
rect 6692 24444 6804 24500
rect 6636 24406 6692 24444
rect 6468 23996 6580 24052
rect 6412 23986 6468 23996
rect 6188 22260 6244 22270
rect 5964 22258 6244 22260
rect 5964 22206 6190 22258
rect 6242 22206 6244 22258
rect 5964 22204 6244 22206
rect 5180 21588 5236 21598
rect 5180 20356 5236 21532
rect 6076 21588 6132 21598
rect 6076 21494 6132 21532
rect 5964 21476 6020 21486
rect 5852 20916 5908 20926
rect 5964 20916 6020 21420
rect 5908 20860 6020 20916
rect 5852 20850 5908 20860
rect 5852 20580 5908 20590
rect 5852 20578 6020 20580
rect 5852 20526 5854 20578
rect 5906 20526 6020 20578
rect 5852 20524 6020 20526
rect 5852 20514 5908 20524
rect 5180 20018 5236 20300
rect 5180 19966 5182 20018
rect 5234 19966 5236 20018
rect 5180 19954 5236 19966
rect 5740 19234 5796 19246
rect 5740 19182 5742 19234
rect 5794 19182 5796 19234
rect 5740 19124 5796 19182
rect 5740 19058 5796 19068
rect 5852 19234 5908 19246
rect 5852 19182 5854 19234
rect 5906 19182 5908 19234
rect 5068 18900 5124 18956
rect 4844 18844 5124 18900
rect 4732 17444 4788 17454
rect 4732 17350 4788 17388
rect 4172 16830 4174 16882
rect 4226 16830 4228 16882
rect 4172 16818 4228 16830
rect 4508 16884 4564 16894
rect 4396 16324 4452 16334
rect 4508 16324 4564 16828
rect 4396 16322 4564 16324
rect 4396 16270 4398 16322
rect 4450 16270 4564 16322
rect 4396 16268 4564 16270
rect 4396 16258 4452 16268
rect 4172 16212 4228 16222
rect 4172 14196 4228 16156
rect 4620 15986 4676 16940
rect 4620 15934 4622 15986
rect 4674 15934 4676 15986
rect 4620 15922 4676 15934
rect 4732 16658 4788 16670
rect 4732 16606 4734 16658
rect 4786 16606 4788 16658
rect 4508 15874 4564 15886
rect 4508 15822 4510 15874
rect 4562 15822 4564 15874
rect 4396 15428 4452 15438
rect 4396 15334 4452 15372
rect 4508 15148 4564 15822
rect 4732 15540 4788 16606
rect 4844 15540 4900 18844
rect 5292 18676 5348 18686
rect 5292 18450 5348 18620
rect 5740 18564 5796 18574
rect 5852 18564 5908 19182
rect 5964 19236 6020 20524
rect 6076 19236 6132 19246
rect 5964 19180 6076 19236
rect 6076 19170 6132 19180
rect 5796 18508 5908 18564
rect 5740 18470 5796 18508
rect 6076 18452 6132 18462
rect 5292 18398 5294 18450
rect 5346 18398 5348 18450
rect 5292 16772 5348 18398
rect 5964 18396 6076 18452
rect 5628 17780 5684 17790
rect 5292 16706 5348 16716
rect 5516 17444 5572 17454
rect 5516 16770 5572 17388
rect 5628 16882 5684 17724
rect 5740 17554 5796 17566
rect 5740 17502 5742 17554
rect 5794 17502 5796 17554
rect 5740 16996 5796 17502
rect 5964 17554 6020 18396
rect 6076 18358 6132 18396
rect 6076 17780 6132 17790
rect 6076 17686 6132 17724
rect 5964 17502 5966 17554
rect 6018 17502 6020 17554
rect 5964 17490 6020 17502
rect 5740 16930 5796 16940
rect 5628 16830 5630 16882
rect 5682 16830 5684 16882
rect 5628 16818 5684 16830
rect 5516 16718 5518 16770
rect 5570 16718 5572 16770
rect 5292 16548 5348 16558
rect 4844 15484 5012 15540
rect 4732 15474 4788 15484
rect 4508 15092 4788 15148
rect 4508 14980 4564 14990
rect 4172 14130 4228 14140
rect 4284 14532 4340 14542
rect 4284 13972 4340 14476
rect 4284 13906 4340 13916
rect 4396 14418 4452 14430
rect 4396 14366 4398 14418
rect 4450 14366 4452 14418
rect 4284 13748 4340 13758
rect 4172 13746 4340 13748
rect 4172 13694 4286 13746
rect 4338 13694 4340 13746
rect 4172 13692 4340 13694
rect 4172 11732 4228 13692
rect 4284 13682 4340 13692
rect 4396 13074 4452 14366
rect 4396 13022 4398 13074
rect 4450 13022 4452 13074
rect 4396 13010 4452 13022
rect 4284 12964 4340 12974
rect 4284 12870 4340 12908
rect 4172 11666 4228 11676
rect 4508 11506 4564 14924
rect 4732 14418 4788 15092
rect 4732 14366 4734 14418
rect 4786 14366 4788 14418
rect 4732 12964 4788 14366
rect 4844 14308 4900 14318
rect 4956 14308 5012 15484
rect 5292 15428 5348 16492
rect 5292 15334 5348 15372
rect 5516 14980 5572 16718
rect 6076 16772 6132 16782
rect 6076 16212 6132 16716
rect 6076 15316 6132 16156
rect 5516 14914 5572 14924
rect 5740 15314 6132 15316
rect 5740 15262 6078 15314
rect 6130 15262 6132 15314
rect 5740 15260 6132 15262
rect 4844 14306 5012 14308
rect 4844 14254 4846 14306
rect 4898 14254 5012 14306
rect 4844 14252 5012 14254
rect 4844 14242 4900 14252
rect 4732 12898 4788 12908
rect 4844 13074 4900 13086
rect 4844 13022 4846 13074
rect 4898 13022 4900 13074
rect 4844 12292 4900 13022
rect 4844 12226 4900 12236
rect 4508 11454 4510 11506
rect 4562 11454 4564 11506
rect 4508 11442 4564 11454
rect 4844 11956 4900 11966
rect 4060 10770 4116 10780
rect 4172 11396 4228 11406
rect 3948 10388 4004 10398
rect 3948 9826 4004 10332
rect 3948 9774 3950 9826
rect 4002 9774 4004 9826
rect 3836 9380 3892 9390
rect 3948 9380 4004 9774
rect 3892 9324 4004 9380
rect 4172 9826 4228 11340
rect 4620 10612 4676 10622
rect 4620 10050 4676 10556
rect 4620 9998 4622 10050
rect 4674 9998 4676 10050
rect 4620 9986 4676 9998
rect 4172 9774 4174 9826
rect 4226 9774 4228 9826
rect 3836 9314 3892 9324
rect 3724 9102 3726 9154
rect 3778 9102 3780 9154
rect 3724 8932 3780 9102
rect 3836 9156 3892 9166
rect 3836 9062 3892 9100
rect 4060 9044 4116 9054
rect 4060 8950 4116 8988
rect 3724 8876 3892 8932
rect 3612 8764 3780 8820
rect 3164 8258 3668 8260
rect 3164 8206 3166 8258
rect 3218 8206 3668 8258
rect 3164 8204 3668 8206
rect 3164 8194 3220 8204
rect 2828 7634 2884 7644
rect 2940 7868 3108 7924
rect 2828 7476 2884 7486
rect 2828 7382 2884 7420
rect 2940 7252 2996 7868
rect 3388 7812 3444 7822
rect 3388 7586 3444 7756
rect 3388 7534 3390 7586
rect 3442 7534 3444 7586
rect 3052 7476 3108 7486
rect 3108 7420 3332 7476
rect 3052 7410 3108 7420
rect 2492 7196 2660 7252
rect 2828 7196 2996 7252
rect 2380 7140 2436 7150
rect 2268 7084 2380 7140
rect 2380 7074 2436 7084
rect 1932 6356 1988 6366
rect 1820 6300 1932 6356
rect 1932 6290 1988 6300
rect 1820 6132 1876 6142
rect 1820 6038 1876 6076
rect 2044 6020 2100 6030
rect 1820 5122 1876 5134
rect 1820 5070 1822 5122
rect 1874 5070 1876 5122
rect 1820 5012 1876 5070
rect 1820 4564 1876 4956
rect 1820 4498 1876 4508
rect 2044 4562 2100 5964
rect 2380 5796 2436 5806
rect 2268 5740 2380 5796
rect 2268 5234 2324 5740
rect 2380 5702 2436 5740
rect 2268 5182 2270 5234
rect 2322 5182 2324 5234
rect 2268 5170 2324 5182
rect 2044 4510 2046 4562
rect 2098 4510 2100 4562
rect 2044 4498 2100 4510
rect 2492 4562 2548 7196
rect 2716 6802 2772 6814
rect 2716 6750 2718 6802
rect 2770 6750 2772 6802
rect 2716 6692 2772 6750
rect 2716 6626 2772 6636
rect 2716 6356 2772 6366
rect 2604 5908 2660 5918
rect 2604 5814 2660 5852
rect 2716 5234 2772 6300
rect 2716 5182 2718 5234
rect 2770 5182 2772 5234
rect 2716 5170 2772 5182
rect 2492 4510 2494 4562
rect 2546 4510 2548 4562
rect 2492 4498 2548 4510
rect 1820 4338 1876 4350
rect 1820 4286 1822 4338
rect 1874 4286 1876 4338
rect 1820 3668 1876 4286
rect 1708 3554 1764 3566
rect 1708 3502 1710 3554
rect 1762 3502 1764 3554
rect 1708 3444 1764 3502
rect 1708 1428 1764 3388
rect 1820 3332 1876 3612
rect 2828 3666 2884 7196
rect 3052 7140 3108 7150
rect 2940 5684 2996 5694
rect 2940 5590 2996 5628
rect 3052 4564 3108 7084
rect 3276 6914 3332 7420
rect 3276 6862 3278 6914
rect 3330 6862 3332 6914
rect 3276 6850 3332 6862
rect 3164 5796 3220 5806
rect 3164 5236 3220 5740
rect 3164 5234 3332 5236
rect 3164 5182 3166 5234
rect 3218 5182 3332 5234
rect 3164 5180 3332 5182
rect 3164 5170 3220 5180
rect 3164 4564 3220 4574
rect 3052 4562 3220 4564
rect 3052 4510 3166 4562
rect 3218 4510 3220 4562
rect 3052 4508 3220 4510
rect 3164 4498 3220 4508
rect 3276 3892 3332 5180
rect 3388 4114 3444 7534
rect 3612 6914 3668 8204
rect 3612 6862 3614 6914
rect 3666 6862 3668 6914
rect 3612 6850 3668 6862
rect 3500 6692 3556 6702
rect 3724 6692 3780 8764
rect 3836 8596 3892 8876
rect 3948 8930 4004 8942
rect 3948 8878 3950 8930
rect 4002 8878 4004 8930
rect 3948 8820 4004 8878
rect 3948 8754 4004 8764
rect 3836 8372 3892 8540
rect 3836 8306 3892 8316
rect 3948 8370 4004 8382
rect 3948 8318 3950 8370
rect 4002 8318 4004 8370
rect 3948 8260 4004 8318
rect 3948 8194 4004 8204
rect 3836 8148 3892 8158
rect 3836 7588 3892 8092
rect 4060 8036 4116 8046
rect 3836 7586 4004 7588
rect 3836 7534 3838 7586
rect 3890 7534 4004 7586
rect 3836 7532 4004 7534
rect 3836 7522 3892 7532
rect 3836 6692 3892 6702
rect 3724 6690 3892 6692
rect 3724 6638 3838 6690
rect 3890 6638 3892 6690
rect 3724 6636 3892 6638
rect 3500 6130 3556 6636
rect 3500 6078 3502 6130
rect 3554 6078 3556 6130
rect 3500 6066 3556 6078
rect 3836 6020 3892 6636
rect 3836 5954 3892 5964
rect 3724 5908 3780 5918
rect 3612 5852 3724 5908
rect 3612 4900 3668 5852
rect 3724 5842 3780 5852
rect 3836 5796 3892 5806
rect 3836 5702 3892 5740
rect 3724 5684 3780 5694
rect 3724 5124 3780 5628
rect 3948 5124 4004 7532
rect 4060 7474 4116 7980
rect 4060 7422 4062 7474
rect 4114 7422 4116 7474
rect 4060 7410 4116 7422
rect 4172 5796 4228 9774
rect 4508 9938 4564 9950
rect 4508 9886 4510 9938
rect 4562 9886 4564 9938
rect 4508 9828 4564 9886
rect 4508 9492 4564 9772
rect 4844 9716 4900 11900
rect 4956 11506 5012 14252
rect 5068 14306 5124 14318
rect 5068 14254 5070 14306
rect 5122 14254 5124 14306
rect 5068 13748 5124 14254
rect 5740 14308 5796 15260
rect 6076 15250 6132 15260
rect 5964 15092 6020 15102
rect 5852 14308 5908 14318
rect 5740 14306 5908 14308
rect 5740 14254 5854 14306
rect 5906 14254 5908 14306
rect 5740 14252 5908 14254
rect 5628 14196 5684 14206
rect 5628 13972 5684 14140
rect 5740 13972 5796 13982
rect 5628 13970 5796 13972
rect 5628 13918 5742 13970
rect 5794 13918 5796 13970
rect 5628 13916 5796 13918
rect 5740 13906 5796 13916
rect 5068 12962 5124 13692
rect 5068 12910 5070 12962
rect 5122 12910 5124 12962
rect 5068 12898 5124 12910
rect 5852 12516 5908 14252
rect 5964 13860 6020 15036
rect 5964 13766 6020 13804
rect 6076 15090 6132 15102
rect 6076 15038 6078 15090
rect 6130 15038 6132 15090
rect 6076 13412 6132 15038
rect 6188 14532 6244 22204
rect 6300 22260 6356 22988
rect 6300 21476 6356 22204
rect 6524 21700 6580 23996
rect 6636 23716 6692 23726
rect 6636 23622 6692 23660
rect 6748 23156 6804 24444
rect 7196 24052 7252 24558
rect 7196 23828 7252 23996
rect 7196 23762 7252 23772
rect 7532 23492 7588 23502
rect 6748 23154 7252 23156
rect 6748 23102 6750 23154
rect 6802 23102 7252 23154
rect 6748 23100 7252 23102
rect 6748 23090 6804 23100
rect 7196 22370 7252 23100
rect 7196 22318 7198 22370
rect 7250 22318 7252 22370
rect 7196 22306 7252 22318
rect 7308 22820 7364 22830
rect 6524 21644 6692 21700
rect 6300 21410 6356 21420
rect 6412 21362 6468 21374
rect 6412 21310 6414 21362
rect 6466 21310 6468 21362
rect 6300 21028 6356 21038
rect 6300 20914 6356 20972
rect 6300 20862 6302 20914
rect 6354 20862 6356 20914
rect 6300 20850 6356 20862
rect 6412 20916 6468 21310
rect 6412 20850 6468 20860
rect 6636 18676 6692 21644
rect 6972 21698 7028 21710
rect 6972 21646 6974 21698
rect 7026 21646 7028 21698
rect 6748 20804 6804 20842
rect 6748 20738 6804 20748
rect 6860 20692 6916 20702
rect 6860 20598 6916 20636
rect 6524 18620 6692 18676
rect 6860 20468 6916 20478
rect 6300 18338 6356 18350
rect 6300 18286 6302 18338
rect 6354 18286 6356 18338
rect 6300 15148 6356 18286
rect 6524 17108 6580 18620
rect 6748 18564 6804 18574
rect 6748 18470 6804 18508
rect 6860 17666 6916 20412
rect 6860 17614 6862 17666
rect 6914 17614 6916 17666
rect 6860 17602 6916 17614
rect 6972 18452 7028 21646
rect 7196 21586 7252 21598
rect 7196 21534 7198 21586
rect 7250 21534 7252 21586
rect 7084 19908 7140 19918
rect 7084 18564 7140 19852
rect 7196 19124 7252 21534
rect 7196 19058 7252 19068
rect 7084 18498 7140 18508
rect 6972 17108 7028 18396
rect 7084 18340 7140 18350
rect 7084 17780 7140 18284
rect 7084 17666 7140 17724
rect 7196 17892 7252 17902
rect 7196 17778 7252 17836
rect 7196 17726 7198 17778
rect 7250 17726 7252 17778
rect 7196 17714 7252 17726
rect 7084 17614 7086 17666
rect 7138 17614 7140 17666
rect 7084 17602 7140 17614
rect 7084 17108 7140 17118
rect 6524 17052 6692 17108
rect 6972 17052 7084 17108
rect 6524 16884 6580 16894
rect 6524 16790 6580 16828
rect 6636 16772 6692 17052
rect 7084 17042 7140 17052
rect 7084 16884 7140 16894
rect 7084 16790 7140 16828
rect 6636 16716 6804 16772
rect 6524 16212 6580 16222
rect 6524 16098 6580 16156
rect 6524 16046 6526 16098
rect 6578 16046 6580 16098
rect 6524 16034 6580 16046
rect 6748 15538 6804 16716
rect 6748 15486 6750 15538
rect 6802 15486 6804 15538
rect 6636 15428 6692 15438
rect 6636 15334 6692 15372
rect 6748 15148 6804 15486
rect 7084 16098 7140 16110
rect 7084 16046 7086 16098
rect 7138 16046 7140 16098
rect 7084 15428 7140 16046
rect 7084 15362 7140 15372
rect 6300 15092 6468 15148
rect 6300 14980 6356 14990
rect 6300 14642 6356 14924
rect 6300 14590 6302 14642
rect 6354 14590 6356 14642
rect 6300 14578 6356 14590
rect 6188 14466 6244 14476
rect 6412 14420 6468 15092
rect 6412 14354 6468 14364
rect 6524 15092 6804 15148
rect 6972 15314 7028 15326
rect 6972 15262 6974 15314
rect 7026 15262 7028 15314
rect 6972 15148 7028 15262
rect 6972 15092 7140 15148
rect 6188 13748 6244 13758
rect 6188 13654 6244 13692
rect 6076 13346 6132 13356
rect 5964 13076 6020 13086
rect 5964 12982 6020 13020
rect 4956 11454 4958 11506
rect 5010 11454 5012 11506
rect 4956 11442 5012 11454
rect 5516 12460 5908 12516
rect 6300 12740 6356 12750
rect 6524 12740 6580 15092
rect 7084 15090 7140 15092
rect 7084 15038 7086 15090
rect 7138 15038 7140 15090
rect 7084 15026 7140 15038
rect 7308 14644 7364 22764
rect 7420 21700 7476 21710
rect 7420 21606 7476 21644
rect 7532 21476 7588 23436
rect 7420 21420 7588 21476
rect 7420 19684 7476 21420
rect 7644 21364 7700 24670
rect 7756 24500 7812 25454
rect 7756 23938 7812 24444
rect 7756 23886 7758 23938
rect 7810 23886 7812 23938
rect 7756 23874 7812 23886
rect 8092 25508 8148 25518
rect 8092 25394 8148 25452
rect 8092 25342 8094 25394
rect 8146 25342 8148 25394
rect 8092 23828 8148 25342
rect 8204 24164 8260 26350
rect 9324 26404 9380 26414
rect 9324 26310 9380 26348
rect 9884 26404 9940 29200
rect 29820 26908 29876 29200
rect 49756 27300 49812 29200
rect 57708 27412 57764 27422
rect 49756 27244 50372 27300
rect 29596 26852 29876 26908
rect 15518 26684 15782 26694
rect 15574 26628 15622 26684
rect 15678 26628 15726 26684
rect 15518 26618 15782 26628
rect 12460 26516 12516 26526
rect 13580 26516 13636 26526
rect 12460 26514 12628 26516
rect 12460 26462 12462 26514
rect 12514 26462 12628 26514
rect 12460 26460 12628 26462
rect 12460 26450 12516 26460
rect 9884 26338 9940 26348
rect 10220 26292 10276 26302
rect 8876 26180 8932 26190
rect 8876 26086 8932 26124
rect 9884 26178 9940 26190
rect 9884 26126 9886 26178
rect 9938 26126 9940 26178
rect 8365 25900 8629 25910
rect 8421 25844 8469 25900
rect 8525 25844 8573 25900
rect 8365 25834 8629 25844
rect 8764 25844 8820 25854
rect 8764 24834 8820 25788
rect 9772 25844 9828 25854
rect 9436 25620 9492 25630
rect 9436 25506 9492 25564
rect 9772 25618 9828 25788
rect 9884 25732 9940 26126
rect 9884 25666 9940 25676
rect 9772 25566 9774 25618
rect 9826 25566 9828 25618
rect 9772 25554 9828 25566
rect 9436 25454 9438 25506
rect 9490 25454 9492 25506
rect 9436 25442 9492 25454
rect 9100 25396 9156 25406
rect 8764 24782 8766 24834
rect 8818 24782 8820 24834
rect 8365 24332 8629 24342
rect 8421 24276 8469 24332
rect 8525 24276 8573 24332
rect 8365 24266 8629 24276
rect 8204 24098 8260 24108
rect 7868 23826 8148 23828
rect 7868 23774 8094 23826
rect 8146 23774 8148 23826
rect 7868 23772 8148 23774
rect 7756 22372 7812 22382
rect 7868 22372 7924 23772
rect 8092 23762 8148 23772
rect 8316 23828 8372 23838
rect 8316 23714 8372 23772
rect 8764 23716 8820 24782
rect 8988 25060 9044 25070
rect 8988 24610 9044 25004
rect 8988 24558 8990 24610
rect 9042 24558 9044 24610
rect 8876 24164 8932 24174
rect 8876 24050 8932 24108
rect 8876 23998 8878 24050
rect 8930 23998 8932 24050
rect 8876 23986 8932 23998
rect 8988 23940 9044 24558
rect 8988 23874 9044 23884
rect 9100 23826 9156 25340
rect 9772 25396 9828 25406
rect 9772 24946 9828 25340
rect 9772 24894 9774 24946
rect 9826 24894 9828 24946
rect 9772 24882 9828 24894
rect 10220 24722 10276 26236
rect 11116 26290 11172 26302
rect 11116 26238 11118 26290
rect 11170 26238 11172 26290
rect 10220 24670 10222 24722
rect 10274 24670 10276 24722
rect 10220 24658 10276 24670
rect 10556 26178 10612 26190
rect 10556 26126 10558 26178
rect 10610 26126 10612 26178
rect 9884 24612 9940 24622
rect 9884 24518 9940 24556
rect 10444 24610 10500 24622
rect 10444 24558 10446 24610
rect 10498 24558 10500 24610
rect 9100 23774 9102 23826
rect 9154 23774 9156 23826
rect 9100 23762 9156 23774
rect 10220 24164 10276 24174
rect 8316 23662 8318 23714
rect 8370 23662 8372 23714
rect 8316 23650 8372 23662
rect 8428 23660 8820 23716
rect 8428 23492 8484 23660
rect 8204 23436 8484 23492
rect 8092 23042 8148 23054
rect 8092 22990 8094 23042
rect 8146 22990 8148 23042
rect 8092 22484 8148 22990
rect 8204 22484 8260 23436
rect 8764 23154 8820 23166
rect 8764 23102 8766 23154
rect 8818 23102 8820 23154
rect 8365 22764 8629 22774
rect 8421 22708 8469 22764
rect 8525 22708 8573 22764
rect 8365 22698 8629 22708
rect 8764 22596 8820 23102
rect 9100 23156 9156 23166
rect 9772 23156 9828 23166
rect 9156 23100 9268 23156
rect 9100 23090 9156 23100
rect 8540 22540 8820 22596
rect 8876 22932 8932 22942
rect 8204 22428 8372 22484
rect 8092 22418 8148 22428
rect 7756 22370 7924 22372
rect 7756 22318 7758 22370
rect 7810 22318 7924 22370
rect 7756 22316 7924 22318
rect 8316 22372 8372 22428
rect 8316 22316 8484 22372
rect 7756 22306 7812 22316
rect 7868 22036 7924 22316
rect 8204 22260 8260 22270
rect 8204 22166 8260 22204
rect 8316 22146 8372 22158
rect 8316 22094 8318 22146
rect 8370 22094 8372 22146
rect 8316 22036 8372 22094
rect 7868 21980 8372 22036
rect 8428 21924 8484 22316
rect 8540 22370 8596 22540
rect 8540 22318 8542 22370
rect 8594 22318 8596 22370
rect 8540 22306 8596 22318
rect 8876 22372 8932 22876
rect 8876 22278 8932 22316
rect 9100 22370 9156 22382
rect 9100 22318 9102 22370
rect 9154 22318 9156 22370
rect 8316 21868 8484 21924
rect 7980 21698 8036 21710
rect 7980 21646 7982 21698
rect 8034 21646 8036 21698
rect 7980 21364 8036 21646
rect 8316 21588 8372 21868
rect 8876 21812 8932 21822
rect 8876 21718 8932 21756
rect 7644 21308 8036 21364
rect 8204 21586 8372 21588
rect 8204 21534 8318 21586
rect 8370 21534 8372 21586
rect 8204 21532 8372 21534
rect 7756 20580 7812 20590
rect 7644 20020 7700 20030
rect 7644 19906 7700 19964
rect 7756 20018 7812 20524
rect 7756 19966 7758 20018
rect 7810 19966 7812 20018
rect 7756 19954 7812 19966
rect 7644 19854 7646 19906
rect 7698 19854 7700 19906
rect 7644 19842 7700 19854
rect 7420 19628 7812 19684
rect 7644 19122 7700 19134
rect 7644 19070 7646 19122
rect 7698 19070 7700 19122
rect 7644 18900 7700 19070
rect 7644 18834 7700 18844
rect 7420 18564 7476 18574
rect 7420 15652 7476 18508
rect 7420 15538 7476 15596
rect 7420 15486 7422 15538
rect 7474 15486 7476 15538
rect 7420 15474 7476 15486
rect 7420 15092 7476 15102
rect 7420 15090 7588 15092
rect 7420 15038 7422 15090
rect 7474 15038 7588 15090
rect 7420 15036 7588 15038
rect 7420 15026 7476 15036
rect 7308 14588 7476 14644
rect 6636 14532 6692 14542
rect 6636 13970 6692 14476
rect 6636 13918 6638 13970
rect 6690 13918 6692 13970
rect 6636 13906 6692 13918
rect 6748 14308 6804 14318
rect 6748 13970 6804 14252
rect 6748 13918 6750 13970
rect 6802 13918 6804 13970
rect 6748 13906 6804 13918
rect 6860 13972 6916 13982
rect 6860 13878 6916 13916
rect 6972 13412 7028 13422
rect 6748 12740 6804 12750
rect 6300 12738 6804 12740
rect 6300 12686 6302 12738
rect 6354 12686 6750 12738
rect 6802 12686 6804 12738
rect 6300 12684 6804 12686
rect 5292 11172 5348 11182
rect 5516 11172 5572 12460
rect 5628 12292 5684 12302
rect 6188 12292 6244 12302
rect 5628 12290 6244 12292
rect 5628 12238 5630 12290
rect 5682 12238 6190 12290
rect 6242 12238 6244 12290
rect 5628 12236 6244 12238
rect 5628 12226 5684 12236
rect 5852 11844 5908 12236
rect 6188 12226 6244 12236
rect 5740 11732 5796 11742
rect 5740 11506 5796 11676
rect 5740 11454 5742 11506
rect 5794 11454 5796 11506
rect 5740 11442 5796 11454
rect 5348 11116 5572 11172
rect 4956 10500 5012 10510
rect 4956 10406 5012 10444
rect 4844 9660 5236 9716
rect 4508 9426 4564 9436
rect 4844 9492 4900 9502
rect 4900 9436 5012 9492
rect 4844 9426 4900 9436
rect 4508 9156 4564 9166
rect 4508 9062 4564 9100
rect 4844 9156 4900 9166
rect 4844 9062 4900 9100
rect 4396 9042 4452 9054
rect 4396 8990 4398 9042
rect 4450 8990 4452 9042
rect 4396 8820 4452 8990
rect 4956 8932 5012 9436
rect 5068 9380 5124 9390
rect 5068 9266 5124 9324
rect 5068 9214 5070 9266
rect 5122 9214 5124 9266
rect 5068 9202 5124 9214
rect 4956 8866 5012 8876
rect 5180 9154 5236 9660
rect 5180 9102 5182 9154
rect 5234 9102 5236 9154
rect 4396 8754 4452 8764
rect 4508 8818 4564 8830
rect 4508 8766 4510 8818
rect 4562 8766 4564 8818
rect 4508 8484 4564 8766
rect 5180 8820 5236 9102
rect 4508 8418 4564 8428
rect 4844 8708 4900 8718
rect 4844 8372 4900 8652
rect 5180 8484 5236 8764
rect 4396 7476 4452 7486
rect 4396 7382 4452 7420
rect 4396 6914 4452 6926
rect 4396 6862 4398 6914
rect 4450 6862 4452 6914
rect 4396 6802 4452 6862
rect 4844 6914 4900 8316
rect 4844 6862 4846 6914
rect 4898 6862 4900 6914
rect 4844 6850 4900 6862
rect 4956 8428 5236 8484
rect 4396 6750 4398 6802
rect 4450 6750 4452 6802
rect 4396 6738 4452 6750
rect 4732 6804 4788 6814
rect 4732 6710 4788 6748
rect 4956 6468 5012 8428
rect 5292 7698 5348 11116
rect 5516 10948 5572 10958
rect 5516 8932 5572 10892
rect 5628 10612 5684 10650
rect 5628 10546 5684 10556
rect 5852 10498 5908 11788
rect 6300 11732 6356 12684
rect 6748 12674 6804 12684
rect 6300 11666 6356 11676
rect 6748 12404 6804 12414
rect 6188 11172 6244 11182
rect 6188 11078 6244 11116
rect 5852 10446 5854 10498
rect 5906 10446 5908 10498
rect 5852 10434 5908 10446
rect 6636 10612 6692 10622
rect 6076 10052 6132 10062
rect 6076 9826 6132 9996
rect 6636 10050 6692 10556
rect 6636 9998 6638 10050
rect 6690 9998 6692 10050
rect 6636 9986 6692 9998
rect 6748 9938 6804 12348
rect 6972 12178 7028 13356
rect 7196 12740 7252 12750
rect 7196 12646 7252 12684
rect 6972 12126 6974 12178
rect 7026 12126 7028 12178
rect 6972 11620 7028 12126
rect 7308 11956 7364 11966
rect 7308 11862 7364 11900
rect 6972 11618 7252 11620
rect 6972 11566 6974 11618
rect 7026 11566 7252 11618
rect 6972 11564 7252 11566
rect 6972 11554 7028 11564
rect 6860 11394 6916 11406
rect 6860 11342 6862 11394
rect 6914 11342 6916 11394
rect 6860 10052 6916 11342
rect 6860 9986 6916 9996
rect 7084 11282 7140 11294
rect 7084 11230 7086 11282
rect 7138 11230 7140 11282
rect 6748 9886 6750 9938
rect 6802 9886 6804 9938
rect 6076 9774 6078 9826
rect 6130 9774 6132 9826
rect 6076 9044 6132 9774
rect 6300 9828 6356 9838
rect 6300 9268 6356 9772
rect 6300 9202 6356 9212
rect 6748 9268 6804 9886
rect 6748 9202 6804 9212
rect 7084 9828 7140 11230
rect 7196 10610 7252 11564
rect 7420 11284 7476 14588
rect 7532 14530 7588 15036
rect 7532 14478 7534 14530
rect 7586 14478 7588 14530
rect 7532 13524 7588 14478
rect 7644 15090 7700 15102
rect 7644 15038 7646 15090
rect 7698 15038 7700 15090
rect 7644 14642 7700 15038
rect 7644 14590 7646 14642
rect 7698 14590 7700 14642
rect 7644 13746 7700 14590
rect 7756 13972 7812 19628
rect 7868 16996 7924 21308
rect 8204 18676 8260 21532
rect 8316 21522 8372 21532
rect 8988 21588 9044 21598
rect 8988 21494 9044 21532
rect 8365 21196 8629 21206
rect 8421 21140 8469 21196
rect 8525 21140 8573 21196
rect 8365 21130 8629 21140
rect 8428 20802 8484 20814
rect 8428 20750 8430 20802
rect 8482 20750 8484 20802
rect 8428 20244 8484 20750
rect 9100 20468 9156 22318
rect 9100 20402 9156 20412
rect 8428 20178 8484 20188
rect 8764 19908 8820 19918
rect 8365 19628 8629 19638
rect 8421 19572 8469 19628
rect 8525 19572 8573 19628
rect 8365 19562 8629 19572
rect 8540 19124 8596 19134
rect 8540 19030 8596 19068
rect 8764 19122 8820 19852
rect 8876 19906 8932 19918
rect 8876 19854 8878 19906
rect 8930 19854 8932 19906
rect 8876 19460 8932 19854
rect 8876 19394 8932 19404
rect 9212 19236 9268 23100
rect 9772 23062 9828 23100
rect 10220 21586 10276 24108
rect 10332 23940 10388 23950
rect 10332 23846 10388 23884
rect 10220 21534 10222 21586
rect 10274 21534 10276 21586
rect 10108 21362 10164 21374
rect 10108 21310 10110 21362
rect 10162 21310 10164 21362
rect 9660 20802 9716 20814
rect 9660 20750 9662 20802
rect 9714 20750 9716 20802
rect 9660 19460 9716 20750
rect 10108 20468 10164 21310
rect 10108 20402 10164 20412
rect 10108 20244 10164 20254
rect 9772 20130 9828 20142
rect 9772 20078 9774 20130
rect 9826 20078 9828 20130
rect 9772 19572 9828 20078
rect 9996 20132 10052 20142
rect 9996 20038 10052 20076
rect 9884 19908 9940 19918
rect 9884 19814 9940 19852
rect 9772 19516 10052 19572
rect 9660 19404 9828 19460
rect 8764 19070 8766 19122
rect 8818 19070 8820 19122
rect 8764 19058 8820 19070
rect 8876 19180 9268 19236
rect 9324 19236 9380 19246
rect 8876 18900 8932 19180
rect 9324 19142 9380 19180
rect 8764 18844 8932 18900
rect 9100 19010 9156 19022
rect 9100 18958 9102 19010
rect 9154 18958 9156 19010
rect 8260 18620 8372 18676
rect 8204 18610 8260 18620
rect 8316 18452 8372 18620
rect 8652 18452 8708 18462
rect 8316 18450 8708 18452
rect 8316 18398 8654 18450
rect 8706 18398 8708 18450
rect 8316 18396 8708 18398
rect 8652 18386 8708 18396
rect 7980 18228 8036 18238
rect 7980 18134 8036 18172
rect 8365 18060 8629 18070
rect 8421 18004 8469 18060
rect 8525 18004 8573 18060
rect 8365 17994 8629 18004
rect 8204 17892 8260 17902
rect 8764 17892 8820 18844
rect 7980 17780 8036 17790
rect 7980 17666 8036 17724
rect 7980 17614 7982 17666
rect 8034 17614 8036 17666
rect 7980 17602 8036 17614
rect 8204 17666 8260 17836
rect 8428 17836 8820 17892
rect 8876 18676 8932 18686
rect 8204 17614 8206 17666
rect 8258 17614 8260 17666
rect 8204 17602 8260 17614
rect 8316 17668 8372 17678
rect 8316 17574 8372 17612
rect 8092 17332 8148 17342
rect 7868 16930 7924 16940
rect 7980 17276 8092 17332
rect 7868 16772 7924 16782
rect 7868 15538 7924 16716
rect 7868 15486 7870 15538
rect 7922 15486 7924 15538
rect 7868 15474 7924 15486
rect 7980 16210 8036 17276
rect 8092 17266 8148 17276
rect 8428 16994 8484 17836
rect 8428 16942 8430 16994
rect 8482 16942 8484 16994
rect 8428 16930 8484 16942
rect 8764 16884 8820 16894
rect 7980 16158 7982 16210
rect 8034 16158 8036 16210
rect 7980 15090 8036 16158
rect 8092 16770 8148 16782
rect 8092 16718 8094 16770
rect 8146 16718 8148 16770
rect 8092 16212 8148 16718
rect 8365 16492 8629 16502
rect 8421 16436 8469 16492
rect 8525 16436 8573 16492
rect 8365 16426 8629 16436
rect 8092 16146 8148 16156
rect 8540 16100 8596 16110
rect 8540 16006 8596 16044
rect 7980 15038 7982 15090
rect 8034 15038 8036 15090
rect 7980 15026 8036 15038
rect 8365 14924 8629 14934
rect 8421 14868 8469 14924
rect 8525 14868 8573 14924
rect 8365 14858 8629 14868
rect 8652 14756 8708 14766
rect 8764 14756 8820 16828
rect 8876 16882 8932 18620
rect 9100 18564 9156 18958
rect 9100 18498 9156 18508
rect 8988 18340 9044 18350
rect 9660 18340 9716 18350
rect 8988 18338 9604 18340
rect 8988 18286 8990 18338
rect 9042 18286 9604 18338
rect 8988 18284 9604 18286
rect 8988 18274 9044 18284
rect 9100 17108 9156 17118
rect 8876 16830 8878 16882
rect 8930 16830 8932 16882
rect 8876 16818 8932 16830
rect 8988 16884 9044 16894
rect 8988 16660 9044 16828
rect 8876 16604 9044 16660
rect 8876 15538 8932 16604
rect 8876 15486 8878 15538
rect 8930 15486 8932 15538
rect 8876 15474 8932 15486
rect 8988 15428 9044 15438
rect 8988 15314 9044 15372
rect 8988 15262 8990 15314
rect 9042 15262 9044 15314
rect 8988 15250 9044 15262
rect 8652 14754 8820 14756
rect 8652 14702 8654 14754
rect 8706 14702 8820 14754
rect 8652 14700 8820 14702
rect 8988 14756 9044 14766
rect 8652 14690 8708 14700
rect 8988 14662 9044 14700
rect 8428 14644 8484 14654
rect 8428 14642 8596 14644
rect 8428 14590 8430 14642
rect 8482 14590 8596 14642
rect 8428 14588 8596 14590
rect 8428 14578 8484 14588
rect 8540 14532 8596 14588
rect 9100 14532 9156 17052
rect 9548 16994 9604 18284
rect 9660 18246 9716 18284
rect 9660 17554 9716 17566
rect 9660 17502 9662 17554
rect 9714 17502 9716 17554
rect 9660 17108 9716 17502
rect 9772 17332 9828 19404
rect 9772 17266 9828 17276
rect 9884 18450 9940 18462
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9660 17052 9828 17108
rect 9548 16942 9550 16994
rect 9602 16942 9604 16994
rect 9548 15314 9604 16942
rect 9660 16884 9716 16894
rect 9660 16790 9716 16828
rect 9772 16772 9828 17052
rect 9772 16706 9828 16716
rect 9660 16098 9716 16110
rect 9660 16046 9662 16098
rect 9714 16046 9716 16098
rect 9660 15428 9716 16046
rect 9660 15362 9716 15372
rect 9548 15262 9550 15314
rect 9602 15262 9604 15314
rect 9548 15250 9604 15262
rect 9884 14756 9940 18398
rect 9996 18228 10052 19516
rect 10108 19234 10164 20188
rect 10220 20020 10276 21534
rect 10332 21474 10388 21486
rect 10332 21422 10334 21474
rect 10386 21422 10388 21474
rect 10332 20580 10388 21422
rect 10332 20130 10388 20524
rect 10332 20078 10334 20130
rect 10386 20078 10388 20130
rect 10332 20066 10388 20078
rect 10220 19954 10276 19964
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 10108 19012 10164 19182
rect 10108 18946 10164 18956
rect 10220 19460 10276 19470
rect 10220 18788 10276 19404
rect 10444 19236 10500 24558
rect 10556 21476 10612 26126
rect 11116 26068 11172 26238
rect 11340 26292 11396 26302
rect 11340 26198 11396 26236
rect 12348 26292 12404 26302
rect 12348 26290 12516 26292
rect 12348 26238 12350 26290
rect 12402 26238 12516 26290
rect 12348 26236 12516 26238
rect 12348 26226 12404 26236
rect 11172 26012 11508 26068
rect 11116 26002 11172 26012
rect 11452 25506 11508 26012
rect 12012 25620 12068 25630
rect 12012 25526 12068 25564
rect 11452 25454 11454 25506
rect 11506 25454 11508 25506
rect 11452 25284 11508 25454
rect 11452 25218 11508 25228
rect 11900 25508 11956 25518
rect 11900 24834 11956 25452
rect 12460 25508 12516 26236
rect 12460 25442 12516 25452
rect 12348 25284 12404 25294
rect 12348 25190 12404 25228
rect 11900 24782 11902 24834
rect 11954 24782 11956 24834
rect 10892 24724 10948 24734
rect 10780 23938 10836 23950
rect 10780 23886 10782 23938
rect 10834 23886 10836 23938
rect 10780 23716 10836 23886
rect 10556 21410 10612 21420
rect 10668 23266 10724 23278
rect 10668 23214 10670 23266
rect 10722 23214 10724 23266
rect 10668 21700 10724 23214
rect 10780 22482 10836 23660
rect 10780 22430 10782 22482
rect 10834 22430 10836 22482
rect 10780 22418 10836 22430
rect 10892 22370 10948 24668
rect 11004 24164 11060 24174
rect 11004 23938 11060 24108
rect 11004 23886 11006 23938
rect 11058 23886 11060 23938
rect 11004 23874 11060 23886
rect 11340 23940 11396 23950
rect 11900 23940 11956 24782
rect 12236 24724 12292 24734
rect 12572 24724 12628 26460
rect 13244 26290 13300 26302
rect 13244 26238 13246 26290
rect 13298 26238 13300 26290
rect 13244 25620 13300 26238
rect 13244 25554 13300 25564
rect 13580 26290 13636 26460
rect 21308 26516 21364 26526
rect 21308 26422 21364 26460
rect 26684 26516 26740 26526
rect 13580 26238 13582 26290
rect 13634 26238 13636 26290
rect 13468 25508 13524 25518
rect 13580 25508 13636 26238
rect 14028 26402 14084 26414
rect 14028 26350 14030 26402
rect 14082 26350 14084 26402
rect 13580 25452 13860 25508
rect 13468 25414 13524 25452
rect 12908 25394 12964 25406
rect 12908 25342 12910 25394
rect 12962 25342 12964 25394
rect 12908 24834 12964 25342
rect 13580 25284 13636 25294
rect 12908 24782 12910 24834
rect 12962 24782 12964 24834
rect 12908 24770 12964 24782
rect 13468 25282 13636 25284
rect 13468 25230 13582 25282
rect 13634 25230 13636 25282
rect 13468 25228 13636 25230
rect 12292 24668 12404 24724
rect 12236 24658 12292 24668
rect 11340 23938 11508 23940
rect 11340 23886 11342 23938
rect 11394 23886 11508 23938
rect 11340 23884 11508 23886
rect 11340 23874 11396 23884
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 22306 10948 22318
rect 11452 23154 11508 23884
rect 11900 23874 11956 23884
rect 12236 24052 12292 24062
rect 12236 23938 12292 23996
rect 12236 23886 12238 23938
rect 12290 23886 12292 23938
rect 12012 23714 12068 23726
rect 12012 23662 12014 23714
rect 12066 23662 12068 23714
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 11452 21924 11508 23102
rect 11676 23380 11732 23390
rect 11676 23042 11732 23324
rect 11676 22990 11678 23042
rect 11730 22990 11732 23042
rect 11676 22978 11732 22990
rect 11900 23156 11956 23166
rect 11900 22596 11956 23100
rect 11452 21858 11508 21868
rect 11564 22594 11956 22596
rect 11564 22542 11902 22594
rect 11954 22542 11956 22594
rect 11564 22540 11956 22542
rect 10668 21586 10724 21644
rect 10668 21534 10670 21586
rect 10722 21534 10724 21586
rect 10556 20020 10612 20030
rect 10556 19926 10612 19964
rect 10444 19170 10500 19180
rect 10556 19124 10612 19134
rect 10668 19124 10724 21534
rect 11564 21588 11620 22540
rect 11900 22530 11956 22540
rect 10780 21476 10836 21486
rect 10836 21420 10948 21476
rect 10780 21410 10836 21420
rect 10892 21028 10948 21420
rect 10556 19122 10724 19124
rect 10556 19070 10558 19122
rect 10610 19070 10724 19122
rect 10556 19068 10724 19070
rect 10780 19794 10836 19806
rect 10780 19742 10782 19794
rect 10834 19742 10836 19794
rect 10556 19058 10612 19068
rect 10780 19012 10836 19742
rect 10220 18450 10276 18732
rect 10220 18398 10222 18450
rect 10274 18398 10276 18450
rect 10220 18386 10276 18398
rect 10332 18900 10388 18910
rect 10332 18564 10388 18844
rect 10780 18676 10836 18956
rect 10780 18610 10836 18620
rect 9996 18172 10164 18228
rect 10108 17556 10164 18172
rect 10220 17668 10276 17678
rect 10332 17668 10388 18508
rect 10668 18228 10724 18238
rect 10668 18134 10724 18172
rect 10220 17666 10388 17668
rect 10220 17614 10222 17666
rect 10274 17614 10388 17666
rect 10220 17612 10388 17614
rect 10444 17666 10500 17678
rect 10444 17614 10446 17666
rect 10498 17614 10500 17666
rect 10220 17602 10276 17612
rect 9996 16324 10052 16334
rect 9996 16210 10052 16268
rect 9996 16158 9998 16210
rect 10050 16158 10052 16210
rect 9996 16146 10052 16158
rect 10108 15538 10164 17500
rect 10444 17444 10500 17614
rect 10444 17378 10500 17388
rect 10892 16772 10948 20972
rect 11452 21474 11508 21486
rect 11452 21422 11454 21474
rect 11506 21422 11508 21474
rect 11004 20690 11060 20702
rect 11004 20638 11006 20690
rect 11058 20638 11060 20690
rect 11004 19458 11060 20638
rect 11452 20244 11508 21422
rect 11564 20802 11620 21532
rect 11676 21924 11732 21934
rect 11676 21364 11732 21868
rect 11900 21700 11956 21710
rect 12012 21700 12068 23662
rect 12236 23604 12292 23886
rect 12348 23826 12404 24668
rect 12572 24658 12628 24668
rect 13356 24724 13412 24734
rect 12908 24052 12964 24062
rect 12908 23958 12964 23996
rect 13356 23940 13412 24668
rect 13356 23874 13412 23884
rect 13468 24612 13524 25228
rect 13580 25218 13636 25228
rect 13468 24276 13524 24556
rect 12348 23774 12350 23826
rect 12402 23774 12404 23826
rect 12348 23762 12404 23774
rect 12236 23538 12292 23548
rect 13132 23268 13188 23278
rect 12684 23156 12740 23166
rect 12684 23062 12740 23100
rect 13020 22146 13076 22158
rect 13020 22094 13022 22146
rect 13074 22094 13076 22146
rect 13020 21924 13076 22094
rect 13020 21858 13076 21868
rect 11900 21698 12068 21700
rect 11900 21646 11902 21698
rect 11954 21646 12068 21698
rect 11900 21644 12068 21646
rect 12796 21810 12852 21822
rect 12796 21758 12798 21810
rect 12850 21758 12852 21810
rect 11900 21634 11956 21644
rect 11788 21586 11844 21598
rect 11788 21534 11790 21586
rect 11842 21534 11844 21586
rect 11788 21476 11844 21534
rect 11900 21476 11956 21486
rect 11788 21420 11900 21476
rect 11900 21410 11956 21420
rect 11676 21308 11844 21364
rect 11564 20750 11566 20802
rect 11618 20750 11620 20802
rect 11564 20738 11620 20750
rect 11452 20178 11508 20188
rect 11004 19406 11006 19458
rect 11058 19406 11060 19458
rect 11004 19394 11060 19406
rect 11228 20020 11284 20030
rect 11116 19236 11172 19246
rect 11004 18340 11060 18350
rect 11004 17780 11060 18284
rect 11004 17686 11060 17724
rect 11004 16996 11060 17006
rect 11004 16902 11060 16940
rect 10892 16436 10948 16716
rect 10892 16212 10948 16380
rect 10668 16210 10948 16212
rect 10668 16158 10894 16210
rect 10946 16158 10948 16210
rect 10668 16156 10948 16158
rect 10108 15486 10110 15538
rect 10162 15486 10164 15538
rect 10108 15474 10164 15486
rect 10556 15652 10612 15662
rect 10556 15426 10612 15596
rect 10556 15374 10558 15426
rect 10610 15374 10612 15426
rect 10556 15362 10612 15374
rect 10668 15314 10724 16156
rect 10892 16146 10948 16156
rect 11116 15988 11172 19180
rect 11228 19234 11284 19964
rect 11788 19460 11844 21308
rect 12796 20802 12852 21758
rect 12796 20750 12798 20802
rect 12850 20750 12852 20802
rect 12796 20738 12852 20750
rect 12796 20578 12852 20590
rect 12796 20526 12798 20578
rect 12850 20526 12852 20578
rect 11228 19182 11230 19234
rect 11282 19182 11284 19234
rect 11228 19170 11284 19182
rect 11452 19404 11844 19460
rect 12572 20018 12628 20030
rect 12572 19966 12574 20018
rect 12626 19966 12628 20018
rect 11452 19122 11508 19404
rect 11452 19070 11454 19122
rect 11506 19070 11508 19122
rect 11452 19058 11508 19070
rect 11788 19236 11844 19246
rect 11564 18450 11620 18462
rect 11564 18398 11566 18450
rect 11618 18398 11620 18450
rect 11228 18338 11284 18350
rect 11228 18286 11230 18338
rect 11282 18286 11284 18338
rect 11228 18116 11284 18286
rect 11564 18340 11620 18398
rect 11564 18274 11620 18284
rect 11284 18060 11508 18116
rect 11228 18050 11284 18060
rect 11228 15988 11284 15998
rect 11116 15986 11284 15988
rect 11116 15934 11230 15986
rect 11282 15934 11284 15986
rect 11116 15932 11284 15934
rect 10668 15262 10670 15314
rect 10722 15262 10724 15314
rect 10668 15148 10724 15262
rect 10332 15092 10724 15148
rect 11004 15652 11060 15662
rect 9884 14690 9940 14700
rect 9996 14868 10052 14878
rect 8540 14476 9156 14532
rect 8092 14418 8148 14430
rect 8092 14366 8094 14418
rect 8146 14366 8148 14418
rect 7756 13916 8036 13972
rect 7644 13694 7646 13746
rect 7698 13694 7700 13746
rect 7644 13682 7700 13694
rect 7868 13746 7924 13758
rect 7868 13694 7870 13746
rect 7922 13694 7924 13746
rect 7868 13524 7924 13694
rect 7532 13468 7924 13524
rect 7980 11732 8036 13916
rect 8092 13636 8148 14366
rect 9548 14418 9604 14430
rect 9548 14366 9550 14418
rect 9602 14366 9604 14418
rect 8092 12740 8148 13580
rect 8204 14308 8260 14318
rect 8204 12962 8260 14252
rect 9212 14306 9268 14318
rect 9212 14254 9214 14306
rect 9266 14254 9268 14306
rect 8988 13748 9044 13758
rect 9212 13748 9268 14254
rect 9436 14308 9492 14318
rect 9436 14214 9492 14252
rect 9548 13970 9604 14366
rect 9548 13918 9550 13970
rect 9602 13918 9604 13970
rect 9548 13906 9604 13918
rect 9772 14196 9828 14206
rect 8988 13746 9268 13748
rect 8988 13694 8990 13746
rect 9042 13694 9268 13746
rect 8988 13692 9268 13694
rect 8988 13682 9044 13692
rect 9660 13636 9716 13646
rect 9660 13542 9716 13580
rect 8764 13524 8820 13534
rect 8764 13430 8820 13468
rect 8365 13356 8629 13366
rect 8421 13300 8469 13356
rect 8525 13300 8573 13356
rect 8365 13290 8629 13300
rect 8204 12910 8206 12962
rect 8258 12910 8260 12962
rect 8204 12898 8260 12910
rect 8316 13074 8372 13086
rect 8316 13022 8318 13074
rect 8370 13022 8372 13074
rect 8316 12740 8372 13022
rect 9436 12852 9492 12862
rect 9436 12758 9492 12796
rect 8092 12684 8372 12740
rect 9660 12404 9716 12414
rect 9660 12310 9716 12348
rect 8988 12180 9044 12190
rect 8092 12068 8148 12078
rect 8092 12066 8260 12068
rect 8092 12014 8094 12066
rect 8146 12014 8260 12066
rect 8092 12012 8260 12014
rect 8092 12002 8148 12012
rect 7980 11676 8148 11732
rect 7868 11394 7924 11406
rect 7868 11342 7870 11394
rect 7922 11342 7924 11394
rect 7420 11228 7812 11284
rect 7196 10558 7198 10610
rect 7250 10558 7252 10610
rect 7196 10546 7252 10558
rect 7420 10612 7476 10622
rect 7420 10518 7476 10556
rect 7756 10276 7812 11228
rect 7868 11060 7924 11342
rect 8092 11172 8148 11676
rect 8204 11396 8260 12012
rect 8540 12066 8596 12078
rect 8540 12014 8542 12066
rect 8594 12014 8596 12066
rect 8540 11956 8596 12014
rect 8988 12066 9044 12124
rect 8988 12014 8990 12066
rect 9042 12014 9044 12066
rect 8540 11900 8820 11956
rect 8764 11844 8820 11900
rect 8365 11788 8629 11798
rect 8421 11732 8469 11788
rect 8525 11732 8573 11788
rect 8365 11722 8629 11732
rect 8204 11330 8260 11340
rect 7868 10994 7924 11004
rect 7980 11116 8148 11172
rect 7756 10220 7924 10276
rect 7756 10052 7812 10062
rect 7084 9154 7140 9772
rect 7644 9826 7700 9838
rect 7644 9774 7646 9826
rect 7698 9774 7700 9826
rect 7084 9102 7086 9154
rect 7138 9102 7140 9154
rect 7084 9090 7140 9102
rect 7532 9268 7588 9278
rect 6076 8978 6132 8988
rect 6524 9044 6580 9054
rect 5740 8932 5796 8942
rect 5516 8930 5796 8932
rect 5516 8878 5742 8930
rect 5794 8878 5796 8930
rect 5516 8876 5796 8878
rect 5292 7646 5294 7698
rect 5346 7646 5348 7698
rect 5292 7634 5348 7646
rect 5404 8596 5460 8606
rect 5404 7476 5460 8540
rect 4732 6412 5012 6468
rect 5068 7420 5460 7476
rect 4732 6130 4788 6412
rect 4732 6078 4734 6130
rect 4786 6078 4788 6130
rect 4732 6066 4788 6078
rect 4844 6132 4900 6142
rect 4172 5730 4228 5740
rect 4732 5346 4788 5358
rect 4732 5294 4734 5346
rect 4786 5294 4788 5346
rect 4172 5124 4228 5134
rect 3948 5122 4228 5124
rect 3948 5070 4174 5122
rect 4226 5070 4228 5122
rect 3948 5068 4228 5070
rect 3724 5058 3780 5068
rect 3612 4844 4004 4900
rect 3388 4062 3390 4114
rect 3442 4062 3444 4114
rect 3388 4050 3444 4062
rect 3612 4226 3668 4238
rect 3612 4174 3614 4226
rect 3666 4174 3668 4226
rect 3612 4114 3668 4174
rect 3612 4062 3614 4114
rect 3666 4062 3668 4114
rect 3612 4050 3668 4062
rect 3276 3836 3556 3892
rect 2828 3614 2830 3666
rect 2882 3614 2884 3666
rect 2828 3602 2884 3614
rect 3500 3666 3556 3836
rect 3500 3614 3502 3666
rect 3554 3614 3556 3666
rect 3500 3602 3556 3614
rect 3948 3666 4004 4844
rect 4172 4788 4228 5068
rect 4172 4722 4228 4732
rect 4620 5124 4676 5134
rect 4396 4564 4452 4574
rect 4396 4470 4452 4508
rect 4620 4338 4676 5068
rect 4620 4286 4622 4338
rect 4674 4286 4676 4338
rect 4620 4274 4676 4286
rect 4732 4340 4788 5294
rect 4844 5348 4900 6076
rect 5068 6130 5124 7420
rect 5516 6692 5572 8876
rect 5740 8866 5796 8876
rect 6524 8820 6580 8988
rect 6412 8818 6580 8820
rect 6412 8766 6526 8818
rect 6578 8766 6580 8818
rect 6412 8764 6580 8766
rect 5740 8372 5796 8382
rect 5740 8278 5796 8316
rect 6300 8260 6356 8270
rect 6300 8146 6356 8204
rect 6412 8258 6468 8764
rect 6524 8754 6580 8764
rect 6636 8932 6692 8942
rect 6412 8206 6414 8258
rect 6466 8206 6468 8258
rect 6412 8194 6468 8206
rect 6300 8094 6302 8146
rect 6354 8094 6356 8146
rect 6076 8036 6132 8046
rect 6300 8036 6356 8094
rect 6636 8036 6692 8876
rect 6860 8818 6916 8830
rect 6860 8766 6862 8818
rect 6914 8766 6916 8818
rect 6860 8596 6916 8766
rect 6860 8530 6916 8540
rect 7420 8260 7476 8270
rect 7420 8166 7476 8204
rect 6748 8148 6804 8158
rect 6748 8054 6804 8092
rect 7308 8148 7364 8158
rect 7308 8054 7364 8092
rect 7532 8036 7588 9212
rect 7644 8818 7700 9774
rect 7756 9714 7812 9996
rect 7756 9662 7758 9714
rect 7810 9662 7812 9714
rect 7756 9650 7812 9662
rect 7644 8766 7646 8818
rect 7698 8766 7700 8818
rect 7644 8596 7700 8766
rect 7644 8530 7700 8540
rect 7756 9156 7812 9166
rect 6076 8034 6244 8036
rect 6076 7982 6078 8034
rect 6130 7982 6244 8034
rect 6076 7980 6244 7982
rect 6300 7980 6692 8036
rect 6076 7970 6132 7980
rect 5628 7924 5684 7934
rect 5628 7698 5684 7868
rect 5628 7646 5630 7698
rect 5682 7646 5684 7698
rect 5628 7634 5684 7646
rect 6188 7700 6244 7980
rect 6188 7644 6580 7700
rect 6188 7476 6244 7486
rect 6244 7420 6468 7476
rect 6188 7382 6244 7420
rect 5516 6626 5572 6636
rect 5740 6692 5796 6702
rect 5068 6078 5070 6130
rect 5122 6078 5124 6130
rect 5068 5682 5124 6078
rect 5516 6132 5572 6142
rect 5516 6038 5572 6076
rect 5740 5908 5796 6636
rect 6412 6690 6468 7420
rect 6524 7362 6580 7644
rect 6524 7310 6526 7362
rect 6578 7310 6580 7362
rect 6524 6802 6580 7310
rect 6524 6750 6526 6802
rect 6578 6750 6580 6802
rect 6524 6738 6580 6750
rect 6412 6638 6414 6690
rect 6466 6638 6468 6690
rect 6412 6626 6468 6638
rect 5740 5842 5796 5852
rect 6188 6578 6244 6590
rect 6188 6526 6190 6578
rect 6242 6526 6244 6578
rect 5068 5630 5070 5682
rect 5122 5630 5124 5682
rect 5068 5618 5124 5630
rect 6076 5794 6132 5806
rect 6076 5742 6078 5794
rect 6130 5742 6132 5794
rect 6076 5682 6132 5742
rect 6076 5630 6078 5682
rect 6130 5630 6132 5682
rect 6076 5618 6132 5630
rect 4844 5292 5236 5348
rect 4844 5122 4900 5292
rect 5068 5124 5124 5134
rect 4844 5070 4846 5122
rect 4898 5070 4900 5122
rect 4844 5058 4900 5070
rect 4956 5068 5068 5124
rect 4956 5010 5012 5068
rect 5068 5058 5124 5068
rect 4956 4958 4958 5010
rect 5010 4958 5012 5010
rect 4956 4946 5012 4958
rect 4956 4788 5012 4798
rect 4956 4562 5012 4732
rect 4956 4510 4958 4562
rect 5010 4510 5012 4562
rect 4956 4498 5012 4510
rect 5180 4564 5236 5292
rect 5740 5124 5796 5134
rect 5180 4470 5236 4508
rect 5292 5122 5796 5124
rect 5292 5070 5742 5122
rect 5794 5070 5796 5122
rect 5292 5068 5796 5070
rect 5292 4562 5348 5068
rect 5740 5058 5796 5068
rect 6188 5124 6244 6526
rect 6636 6130 6692 7980
rect 7420 7980 7588 8036
rect 7644 8034 7700 8046
rect 7644 7982 7646 8034
rect 7698 7982 7700 8034
rect 7084 7476 7140 7486
rect 7084 7474 7252 7476
rect 7084 7422 7086 7474
rect 7138 7422 7252 7474
rect 7084 7420 7252 7422
rect 7084 7410 7140 7420
rect 7196 7250 7252 7420
rect 7196 7198 7198 7250
rect 7250 7198 7252 7250
rect 7196 7186 7252 7198
rect 7420 6692 7476 7980
rect 7532 7812 7588 7822
rect 7532 7698 7588 7756
rect 7532 7646 7534 7698
rect 7586 7646 7588 7698
rect 7532 7634 7588 7646
rect 6636 6078 6638 6130
rect 6690 6078 6692 6130
rect 6636 6066 6692 6078
rect 6972 6580 7028 6590
rect 6972 6130 7028 6524
rect 7420 6468 7476 6636
rect 7532 6692 7588 6702
rect 7644 6692 7700 7982
rect 7756 8034 7812 9100
rect 7756 7982 7758 8034
rect 7810 7982 7812 8034
rect 7756 7812 7812 7982
rect 7756 7746 7812 7756
rect 7868 7700 7924 10220
rect 7980 9266 8036 11116
rect 8316 10836 8372 10846
rect 8204 10612 8260 10622
rect 8092 9604 8148 9614
rect 8092 9510 8148 9548
rect 7980 9214 7982 9266
rect 8034 9214 8036 9266
rect 7980 9202 8036 9214
rect 8204 9044 8260 10556
rect 8316 10386 8372 10780
rect 8316 10334 8318 10386
rect 8370 10334 8372 10386
rect 8316 10322 8372 10334
rect 8365 10220 8629 10230
rect 8421 10164 8469 10220
rect 8525 10164 8573 10220
rect 8365 10154 8629 10164
rect 8764 9716 8820 11788
rect 8876 9716 8932 9726
rect 8764 9714 8932 9716
rect 8764 9662 8878 9714
rect 8930 9662 8932 9714
rect 8764 9660 8932 9662
rect 7980 8988 8260 9044
rect 7980 8258 8036 8988
rect 8540 8932 8596 8942
rect 8876 8932 8932 9660
rect 8988 9156 9044 12014
rect 9548 12068 9604 12078
rect 9436 11396 9492 11406
rect 9436 11302 9492 11340
rect 9100 11282 9156 11294
rect 9100 11230 9102 11282
rect 9154 11230 9156 11282
rect 9100 10052 9156 11230
rect 9100 9986 9156 9996
rect 9436 10052 9492 10062
rect 9548 10052 9604 12012
rect 9660 11844 9716 11854
rect 9660 11618 9716 11788
rect 9660 11566 9662 11618
rect 9714 11566 9716 11618
rect 9660 11554 9716 11566
rect 9772 11620 9828 14140
rect 9884 13076 9940 13086
rect 9996 13076 10052 14812
rect 10332 13748 10388 15092
rect 11004 14644 11060 15596
rect 11228 15148 11284 15932
rect 11452 15314 11508 18060
rect 11788 17668 11844 19180
rect 12012 19124 12068 19134
rect 11900 18450 11956 18462
rect 11900 18398 11902 18450
rect 11954 18398 11956 18450
rect 11900 17892 11956 18398
rect 11900 17826 11956 17836
rect 12012 18340 12068 19068
rect 12012 17778 12068 18284
rect 12460 18564 12516 18574
rect 12012 17726 12014 17778
rect 12066 17726 12068 17778
rect 12012 17714 12068 17726
rect 12348 18228 12404 18238
rect 11788 17602 11844 17612
rect 12348 17666 12404 18172
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 11676 17444 11732 17454
rect 11452 15262 11454 15314
rect 11506 15262 11508 15314
rect 11228 15092 11396 15148
rect 10780 14530 10836 14542
rect 10780 14478 10782 14530
rect 10834 14478 10836 14530
rect 10444 14308 10500 14318
rect 10444 14306 10612 14308
rect 10444 14254 10446 14306
rect 10498 14254 10612 14306
rect 10444 14252 10612 14254
rect 10444 14242 10500 14252
rect 10444 13748 10500 13758
rect 10332 13746 10500 13748
rect 10332 13694 10446 13746
rect 10498 13694 10500 13746
rect 10332 13692 10500 13694
rect 10332 13522 10388 13534
rect 10332 13470 10334 13522
rect 10386 13470 10388 13522
rect 10332 13412 10388 13470
rect 9884 13074 10052 13076
rect 9884 13022 9886 13074
rect 9938 13022 10052 13074
rect 9884 13020 10052 13022
rect 10220 13356 10388 13412
rect 9884 13010 9940 13020
rect 10108 12066 10164 12078
rect 10108 12014 10110 12066
rect 10162 12014 10164 12066
rect 10108 11844 10164 12014
rect 10108 11778 10164 11788
rect 9772 11554 9828 11564
rect 9996 11172 10052 11182
rect 9996 11170 10164 11172
rect 9996 11118 9998 11170
rect 10050 11118 10164 11170
rect 9996 11116 10164 11118
rect 9996 11106 10052 11116
rect 9436 10050 9604 10052
rect 9436 9998 9438 10050
rect 9490 9998 9604 10050
rect 9436 9996 9604 9998
rect 9436 9986 9492 9996
rect 8988 9090 9044 9100
rect 9100 9828 9156 9838
rect 8596 8876 8932 8932
rect 8988 8932 9044 8942
rect 9100 8932 9156 9772
rect 8988 8930 9156 8932
rect 8988 8878 8990 8930
rect 9042 8878 9156 8930
rect 8988 8876 9156 8878
rect 8540 8838 8596 8876
rect 8988 8818 9044 8876
rect 8988 8766 8990 8818
rect 9042 8766 9044 8818
rect 8988 8754 9044 8766
rect 8365 8652 8629 8662
rect 8421 8596 8469 8652
rect 8525 8596 8573 8652
rect 8365 8586 8629 8596
rect 8876 8596 8932 8606
rect 7980 8206 7982 8258
rect 8034 8206 8036 8258
rect 7980 8148 8036 8206
rect 8204 8260 8260 8270
rect 8204 8166 8260 8204
rect 7980 8082 8036 8092
rect 8876 8146 8932 8540
rect 9436 8258 9492 8270
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 8876 8094 8878 8146
rect 8930 8094 8932 8146
rect 8876 8082 8932 8094
rect 9212 8148 9268 8158
rect 9212 8054 9268 8092
rect 7980 7700 8036 7710
rect 7868 7698 8036 7700
rect 7868 7646 7982 7698
rect 8034 7646 8036 7698
rect 7868 7644 8036 7646
rect 7980 7634 8036 7644
rect 8428 7700 8484 7710
rect 8428 7606 8484 7644
rect 9436 7698 9492 8206
rect 9436 7646 9438 7698
rect 9490 7646 9492 7698
rect 9436 7634 9492 7646
rect 9548 7476 9604 9996
rect 9660 10948 9716 10958
rect 9660 10722 9716 10892
rect 9660 10670 9662 10722
rect 9714 10670 9716 10722
rect 9660 9268 9716 10670
rect 10108 10612 10164 11116
rect 9884 10386 9940 10398
rect 9884 10334 9886 10386
rect 9938 10334 9940 10386
rect 9884 9828 9940 10334
rect 9996 9828 10052 9838
rect 9940 9826 10052 9828
rect 9940 9774 9998 9826
rect 10050 9774 10052 9826
rect 9940 9772 10052 9774
rect 9884 9762 9940 9772
rect 9996 9762 10052 9772
rect 10108 9492 10164 10556
rect 9660 9174 9716 9212
rect 9772 9380 9828 9390
rect 9772 8708 9828 9324
rect 10108 9266 10164 9436
rect 10108 9214 10110 9266
rect 10162 9214 10164 9266
rect 10108 9202 10164 9214
rect 10220 10388 10276 13356
rect 10332 13076 10388 13086
rect 10332 12982 10388 13020
rect 10444 12404 10500 13692
rect 10444 12338 10500 12348
rect 10556 13636 10612 14252
rect 10780 13860 10836 14478
rect 10780 13794 10836 13804
rect 11004 14530 11060 14588
rect 11004 14478 11006 14530
rect 11058 14478 11060 14530
rect 10668 13636 10724 13646
rect 10556 13580 10668 13636
rect 10556 12402 10612 13580
rect 10668 13542 10724 13580
rect 10780 13522 10836 13534
rect 10780 13470 10782 13522
rect 10834 13470 10836 13522
rect 10780 13412 10836 13470
rect 10780 13346 10836 13356
rect 11004 12962 11060 14478
rect 11340 14532 11396 15092
rect 11452 14868 11508 15262
rect 11564 15538 11620 15550
rect 11564 15486 11566 15538
rect 11618 15486 11620 15538
rect 11564 15316 11620 15486
rect 11676 15540 11732 17388
rect 12348 17332 12404 17614
rect 12348 17266 12404 17276
rect 12012 16994 12068 17006
rect 12012 16942 12014 16994
rect 12066 16942 12068 16994
rect 11676 15484 11844 15540
rect 11676 15316 11732 15326
rect 11564 15260 11676 15316
rect 11452 14802 11508 14812
rect 11452 14532 11508 14542
rect 11340 14530 11452 14532
rect 11340 14478 11342 14530
rect 11394 14478 11452 14530
rect 11340 14476 11452 14478
rect 11340 14466 11396 14476
rect 11116 14306 11172 14318
rect 11116 14254 11118 14306
rect 11170 14254 11172 14306
rect 11116 13746 11172 14254
rect 11116 13694 11118 13746
rect 11170 13694 11172 13746
rect 11116 13682 11172 13694
rect 11340 13746 11396 13758
rect 11340 13694 11342 13746
rect 11394 13694 11396 13746
rect 11340 13412 11396 13694
rect 11340 13346 11396 13356
rect 11116 13076 11172 13086
rect 11116 12982 11172 13020
rect 11004 12910 11006 12962
rect 11058 12910 11060 12962
rect 10556 12350 10558 12402
rect 10610 12350 10612 12402
rect 10556 12338 10612 12350
rect 10668 12850 10724 12862
rect 10668 12798 10670 12850
rect 10722 12798 10724 12850
rect 10668 12180 10724 12798
rect 11004 12628 11060 12910
rect 11340 12964 11396 12974
rect 11452 12964 11508 14476
rect 11564 14530 11620 14542
rect 11564 14478 11566 14530
rect 11618 14478 11620 14530
rect 11564 14420 11620 14478
rect 11564 14354 11620 14364
rect 11676 13746 11732 15260
rect 11788 15148 11844 15484
rect 12012 15428 12068 16942
rect 12348 16100 12404 16110
rect 12348 16006 12404 16044
rect 12012 15362 12068 15372
rect 12348 15316 12404 15326
rect 12348 15222 12404 15260
rect 11788 15092 12292 15148
rect 12124 14642 12180 14654
rect 12124 14590 12126 14642
rect 12178 14590 12180 14642
rect 12124 14532 12180 14590
rect 12124 14466 12180 14476
rect 12236 14530 12292 15092
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 12236 14196 12292 14478
rect 11676 13694 11678 13746
rect 11730 13694 11732 13746
rect 11676 13682 11732 13694
rect 12124 14140 12292 14196
rect 12124 13636 12180 14140
rect 12460 14084 12516 18508
rect 11340 12962 11508 12964
rect 11340 12910 11342 12962
rect 11394 12910 11508 12962
rect 11340 12908 11508 12910
rect 11676 12962 11732 12974
rect 11676 12910 11678 12962
rect 11730 12910 11732 12962
rect 11340 12898 11396 12908
rect 11004 12572 11508 12628
rect 11004 12404 11060 12414
rect 10668 12114 10724 12124
rect 10780 12348 11004 12404
rect 10780 11506 10836 12348
rect 11004 12310 11060 12348
rect 10780 11454 10782 11506
rect 10834 11454 10836 11506
rect 10780 11442 10836 11454
rect 11228 11506 11284 12572
rect 11452 12402 11508 12572
rect 11452 12350 11454 12402
rect 11506 12350 11508 12402
rect 11452 12338 11508 12350
rect 11676 12404 11732 12910
rect 12124 12964 12180 13580
rect 12236 14028 12516 14084
rect 12236 13186 12292 14028
rect 12348 13860 12404 13870
rect 12572 13860 12628 19966
rect 12796 20020 12852 20526
rect 12796 19954 12852 19964
rect 12908 20018 12964 20030
rect 12908 19966 12910 20018
rect 12962 19966 12964 20018
rect 12908 18340 12964 19966
rect 12684 18284 12964 18340
rect 12684 17106 12740 18284
rect 12908 17668 12964 17678
rect 12908 17574 12964 17612
rect 13020 17220 13076 17230
rect 12684 17054 12686 17106
rect 12738 17054 12740 17106
rect 12684 17042 12740 17054
rect 12908 17108 12964 17118
rect 12684 16882 12740 16894
rect 12684 16830 12686 16882
rect 12738 16830 12740 16882
rect 12684 15986 12740 16830
rect 12684 15934 12686 15986
rect 12738 15934 12740 15986
rect 12684 15316 12740 15934
rect 12684 15250 12740 15260
rect 12908 14418 12964 17052
rect 12908 14366 12910 14418
rect 12962 14366 12964 14418
rect 12908 14354 12964 14366
rect 12348 13858 12628 13860
rect 12348 13806 12350 13858
rect 12402 13806 12628 13858
rect 12348 13804 12628 13806
rect 12348 13794 12404 13804
rect 12236 13134 12238 13186
rect 12290 13134 12292 13186
rect 12236 13122 12292 13134
rect 12684 13746 12740 13758
rect 12684 13694 12686 13746
rect 12738 13694 12740 13746
rect 12684 13076 12740 13694
rect 12684 13010 12740 13020
rect 12796 13634 12852 13646
rect 12796 13582 12798 13634
rect 12850 13582 12852 13634
rect 12236 12964 12292 12974
rect 12124 12962 12292 12964
rect 12124 12910 12238 12962
rect 12290 12910 12292 12962
rect 12124 12908 12292 12910
rect 12236 12852 12292 12908
rect 12572 12962 12628 12974
rect 12572 12910 12574 12962
rect 12626 12910 12628 12962
rect 12236 12796 12516 12852
rect 11676 12338 11732 12348
rect 12236 12404 12292 12414
rect 12236 12178 12292 12348
rect 12236 12126 12238 12178
rect 12290 12126 12292 12178
rect 12236 12114 12292 12126
rect 12460 12180 12516 12796
rect 12572 12404 12628 12910
rect 12572 12348 12740 12404
rect 12572 12180 12628 12190
rect 12460 12178 12628 12180
rect 12460 12126 12574 12178
rect 12626 12126 12628 12178
rect 12460 12124 12628 12126
rect 12012 12066 12068 12078
rect 12012 12014 12014 12066
rect 12066 12014 12068 12066
rect 11228 11454 11230 11506
rect 11282 11454 11284 11506
rect 11228 11442 11284 11454
rect 11340 11620 11396 11630
rect 10668 10612 10724 10622
rect 10668 10610 10948 10612
rect 10668 10558 10670 10610
rect 10722 10558 10948 10610
rect 10668 10556 10948 10558
rect 9996 9044 10052 9054
rect 9996 8950 10052 8988
rect 9660 8652 9828 8708
rect 9660 8596 9716 8652
rect 9660 7698 9716 8540
rect 9772 8260 9828 8270
rect 9772 8166 9828 8204
rect 10220 8036 10276 10332
rect 10556 10500 10612 10510
rect 10444 9828 10500 9838
rect 10444 9734 10500 9772
rect 10220 7970 10276 7980
rect 10332 9042 10388 9054
rect 10332 8990 10334 9042
rect 10386 8990 10388 9042
rect 10332 8370 10388 8990
rect 10332 8318 10334 8370
rect 10386 8318 10388 8370
rect 9660 7646 9662 7698
rect 9714 7646 9716 7698
rect 9660 7634 9716 7646
rect 9772 7476 9828 7486
rect 9548 7474 10052 7476
rect 9548 7422 9774 7474
rect 9826 7422 10052 7474
rect 9548 7420 10052 7422
rect 9772 7410 9828 7420
rect 7756 7250 7812 7262
rect 7756 7198 7758 7250
rect 7810 7198 7812 7250
rect 7756 6802 7812 7198
rect 8365 7084 8629 7094
rect 8421 7028 8469 7084
rect 8525 7028 8573 7084
rect 8365 7018 8629 7028
rect 7756 6750 7758 6802
rect 7810 6750 7812 6802
rect 7756 6738 7812 6750
rect 9996 6802 10052 7420
rect 10332 7474 10388 8318
rect 10556 8372 10612 10444
rect 10668 9380 10724 10556
rect 10892 10500 10948 10556
rect 11228 10610 11284 10622
rect 11228 10558 11230 10610
rect 11282 10558 11284 10610
rect 11228 10500 11284 10558
rect 10892 10444 11284 10500
rect 10780 10386 10836 10398
rect 11340 10388 11396 11564
rect 11788 11620 11844 11630
rect 11788 11526 11844 11564
rect 10780 10334 10782 10386
rect 10834 10334 10836 10386
rect 10780 9492 10836 10334
rect 11228 10332 11396 10388
rect 11452 11394 11508 11406
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11228 9714 11284 10332
rect 11228 9662 11230 9714
rect 11282 9662 11284 9714
rect 11228 9650 11284 9662
rect 11452 9492 11508 11342
rect 11676 11172 11732 11182
rect 11676 11078 11732 11116
rect 11788 10724 11844 10734
rect 11788 10052 11844 10668
rect 10780 9436 11508 9492
rect 11564 9996 11844 10052
rect 12012 10612 12068 12014
rect 12124 11844 12180 11854
rect 12124 10724 12180 11788
rect 12572 11508 12628 12124
rect 12684 11844 12740 12348
rect 12796 12402 12852 13582
rect 13020 12404 13076 17164
rect 12796 12350 12798 12402
rect 12850 12350 12852 12402
rect 12796 12338 12852 12350
rect 12908 12348 13076 12404
rect 12684 11778 12740 11788
rect 12908 11620 12964 12348
rect 12908 11554 12964 11564
rect 12572 11414 12628 11452
rect 13020 11508 13076 11518
rect 13020 11414 13076 11452
rect 12124 10630 12180 10668
rect 12572 10724 12628 10734
rect 12572 10630 12628 10668
rect 11564 9938 11620 9996
rect 11564 9886 11566 9938
rect 11618 9886 11620 9938
rect 10668 9314 10724 9324
rect 10668 9156 10724 9166
rect 10668 9062 10724 9100
rect 11228 9156 11284 9166
rect 11228 9062 11284 9100
rect 10780 9044 10836 9054
rect 10780 9042 10948 9044
rect 10780 8990 10782 9042
rect 10834 8990 10948 9042
rect 10780 8988 10948 8990
rect 10780 8978 10836 8988
rect 10556 8306 10612 8316
rect 10668 8818 10724 8830
rect 10668 8766 10670 8818
rect 10722 8766 10724 8818
rect 10332 7422 10334 7474
rect 10386 7422 10388 7474
rect 10332 7410 10388 7422
rect 10444 8260 10500 8270
rect 10444 7476 10500 8204
rect 10556 8148 10612 8158
rect 10668 8148 10724 8766
rect 10612 8092 10724 8148
rect 10780 8482 10836 8494
rect 10780 8430 10782 8482
rect 10834 8430 10836 8482
rect 10556 8082 10612 8092
rect 10556 7476 10612 7486
rect 10444 7474 10612 7476
rect 10444 7422 10558 7474
rect 10610 7422 10612 7474
rect 10444 7420 10612 7422
rect 10556 7410 10612 7420
rect 9996 6750 9998 6802
rect 10050 6750 10052 6802
rect 7532 6690 7700 6692
rect 7532 6638 7534 6690
rect 7586 6638 7700 6690
rect 7532 6636 7700 6638
rect 7532 6626 7588 6636
rect 7420 6412 7812 6468
rect 6972 6078 6974 6130
rect 7026 6078 7028 6130
rect 6972 6066 7028 6078
rect 7756 6130 7812 6412
rect 7756 6078 7758 6130
rect 7810 6078 7812 6130
rect 7756 5908 7812 6078
rect 7756 5842 7812 5852
rect 7868 6466 7924 6478
rect 7868 6414 7870 6466
rect 7922 6414 7924 6466
rect 7868 5796 7924 6414
rect 8428 6132 8484 6142
rect 7868 5730 7924 5740
rect 7980 6130 8484 6132
rect 7980 6078 8430 6130
rect 8482 6078 8484 6130
rect 7980 6076 8484 6078
rect 7308 5236 7364 5246
rect 7308 5142 7364 5180
rect 6188 5030 6244 5068
rect 6636 5012 6692 5022
rect 6076 4788 6132 4798
rect 5292 4510 5294 4562
rect 5346 4510 5348 4562
rect 5292 4498 5348 4510
rect 5628 4564 5684 4574
rect 5628 4470 5684 4508
rect 6076 4564 6132 4732
rect 6076 4508 6580 4564
rect 4732 4274 4788 4284
rect 6076 4338 6132 4508
rect 6076 4286 6078 4338
rect 6130 4286 6132 4338
rect 6076 4274 6132 4286
rect 6300 4340 6356 4350
rect 4060 4226 4116 4238
rect 4060 4174 4062 4226
rect 4114 4174 4116 4226
rect 4060 4114 4116 4174
rect 4060 4062 4062 4114
rect 4114 4062 4116 4114
rect 4060 4050 4116 4062
rect 3948 3614 3950 3666
rect 4002 3614 4004 3666
rect 3948 3602 4004 3614
rect 4732 3668 4788 3678
rect 4732 3574 4788 3612
rect 6300 3554 6356 4284
rect 6300 3502 6302 3554
rect 6354 3502 6356 3554
rect 6300 3490 6356 3502
rect 6524 3554 6580 4508
rect 6636 4562 6692 4956
rect 6636 4510 6638 4562
rect 6690 4510 6692 4562
rect 6636 4498 6692 4510
rect 7196 4564 7252 4574
rect 6860 4340 6916 4350
rect 6860 3778 6916 4284
rect 6860 3726 6862 3778
rect 6914 3726 6916 3778
rect 6860 3714 6916 3726
rect 7196 3668 7252 4508
rect 7532 4340 7588 4350
rect 7532 4246 7588 4284
rect 7980 4338 8036 6076
rect 8428 6066 8484 6076
rect 9996 6132 10052 6750
rect 10780 6132 10836 8430
rect 10892 8036 10948 8988
rect 11228 8370 11284 8382
rect 11228 8318 11230 8370
rect 11282 8318 11284 8370
rect 11228 8148 11284 8318
rect 11340 8258 11396 9436
rect 11340 8206 11342 8258
rect 11394 8206 11396 8258
rect 11340 8194 11396 8206
rect 11564 8260 11620 9886
rect 12012 9044 12068 10556
rect 13020 10610 13076 10622
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 12796 10386 12852 10398
rect 12796 10334 12798 10386
rect 12850 10334 12852 10386
rect 12796 9940 12852 10334
rect 13020 10388 13076 10558
rect 13020 10322 13076 10332
rect 12796 9874 12852 9884
rect 12572 9602 12628 9614
rect 12572 9550 12574 9602
rect 12626 9550 12628 9602
rect 12572 9156 12628 9550
rect 12572 9090 12628 9100
rect 12012 8978 12068 8988
rect 12908 8820 12964 8830
rect 12908 8370 12964 8764
rect 12908 8318 12910 8370
rect 12962 8318 12964 8370
rect 12908 8306 12964 8318
rect 11564 8194 11620 8204
rect 12460 8260 12516 8270
rect 12460 8166 12516 8204
rect 11228 8082 11284 8092
rect 10892 7970 10948 7980
rect 13132 7924 13188 23212
rect 13468 23266 13524 24220
rect 13468 23214 13470 23266
rect 13522 23214 13524 23266
rect 13468 23202 13524 23214
rect 13580 23714 13636 23726
rect 13580 23662 13582 23714
rect 13634 23662 13636 23714
rect 13580 23604 13636 23662
rect 13580 22372 13636 23548
rect 13468 22370 13636 22372
rect 13468 22318 13582 22370
rect 13634 22318 13636 22370
rect 13468 22316 13636 22318
rect 13468 22260 13524 22316
rect 13580 22306 13636 22316
rect 13692 22372 13748 22382
rect 13468 22194 13524 22204
rect 13692 22258 13748 22316
rect 13692 22206 13694 22258
rect 13746 22206 13748 22258
rect 13692 22148 13748 22206
rect 13692 22082 13748 22092
rect 13804 22146 13860 25452
rect 14028 24722 14084 26350
rect 16044 26404 16100 26414
rect 15036 26068 15092 26078
rect 15036 25974 15092 26012
rect 14364 25620 14420 25630
rect 14364 25506 14420 25564
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 14476 25508 14532 25518
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 13804 22094 13806 22146
rect 13858 22094 13860 22146
rect 13804 22082 13860 22094
rect 13916 24610 13972 24622
rect 13916 24558 13918 24610
rect 13970 24558 13972 24610
rect 13804 21924 13860 21934
rect 13804 21700 13860 21868
rect 13692 18452 13748 18462
rect 13692 18358 13748 18396
rect 13468 16436 13524 16446
rect 13356 16100 13412 16110
rect 13356 15148 13412 16044
rect 13468 16098 13524 16380
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 13468 16034 13524 16046
rect 13580 15988 13636 15998
rect 13356 15092 13524 15148
rect 13468 14644 13524 15092
rect 13468 14578 13524 14588
rect 13580 14642 13636 15932
rect 13804 15148 13860 21644
rect 13916 21588 13972 24558
rect 14028 24164 14084 24670
rect 14084 24108 14308 24164
rect 14028 24098 14084 24108
rect 13916 21494 13972 21532
rect 14028 23940 14084 23950
rect 14028 20802 14084 23884
rect 14028 20750 14030 20802
rect 14082 20750 14084 20802
rect 14028 20738 14084 20750
rect 14140 22596 14196 22606
rect 14140 18676 14196 22540
rect 14252 22260 14308 24108
rect 14476 23940 14532 25452
rect 15148 25508 15204 25518
rect 15148 25414 15204 25452
rect 15518 25116 15782 25126
rect 15574 25060 15622 25116
rect 15678 25060 15726 25116
rect 15518 25050 15782 25060
rect 14924 24724 14980 24734
rect 15148 24724 15204 24734
rect 14924 24722 15092 24724
rect 14924 24670 14926 24722
rect 14978 24670 15092 24722
rect 14924 24668 15092 24670
rect 14924 24658 14980 24668
rect 14476 23874 14532 23884
rect 14588 24610 14644 24622
rect 14588 24558 14590 24610
rect 14642 24558 14644 24610
rect 14476 23154 14532 23166
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 14252 22258 14420 22260
rect 14252 22206 14254 22258
rect 14306 22206 14420 22258
rect 14252 22204 14420 22206
rect 14252 22194 14308 22204
rect 14364 21698 14420 22204
rect 14476 21812 14532 23102
rect 14476 21746 14532 21756
rect 14364 21646 14366 21698
rect 14418 21646 14420 21698
rect 14364 21634 14420 21646
rect 14588 20690 14644 24558
rect 14924 23938 14980 23950
rect 14924 23886 14926 23938
rect 14978 23886 14980 23938
rect 14924 22148 14980 23886
rect 15036 22596 15092 24668
rect 15148 24630 15204 24668
rect 16044 24724 16100 26348
rect 16380 26404 16436 26414
rect 16380 26310 16436 26348
rect 20748 26404 20804 26414
rect 20748 26310 20804 26348
rect 21532 26404 21588 26414
rect 16268 26292 16324 26302
rect 16268 25396 16324 26236
rect 17500 26292 17556 26302
rect 17164 25508 17220 25518
rect 17164 25506 17444 25508
rect 17164 25454 17166 25506
rect 17218 25454 17444 25506
rect 17164 25452 17444 25454
rect 17164 25442 17220 25452
rect 16268 25330 16324 25340
rect 16716 25396 16772 25406
rect 16716 25302 16772 25340
rect 16492 25284 16548 25294
rect 16492 25190 16548 25228
rect 16604 25282 16660 25294
rect 16604 25230 16606 25282
rect 16658 25230 16660 25282
rect 16044 24658 16100 24668
rect 16156 24610 16212 24622
rect 16156 24558 16158 24610
rect 16210 24558 16212 24610
rect 15708 24500 15764 24510
rect 15260 24050 15316 24062
rect 15260 23998 15262 24050
rect 15314 23998 15316 24050
rect 15260 23716 15316 23998
rect 15708 23938 15764 24444
rect 16156 24388 16212 24558
rect 15708 23886 15710 23938
rect 15762 23886 15764 23938
rect 15708 23874 15764 23886
rect 16044 24332 16212 24388
rect 15260 23650 15316 23660
rect 16044 23828 16100 24332
rect 16156 24164 16212 24174
rect 16156 23940 16212 24108
rect 16156 23938 16324 23940
rect 16156 23886 16158 23938
rect 16210 23886 16324 23938
rect 16156 23884 16324 23886
rect 16156 23874 16212 23884
rect 15518 23548 15782 23558
rect 15574 23492 15622 23548
rect 15678 23492 15726 23548
rect 15518 23482 15782 23492
rect 15036 22484 15092 22540
rect 16044 22596 16100 23772
rect 16044 22530 16100 22540
rect 16156 23266 16212 23278
rect 16156 23214 16158 23266
rect 16210 23214 16212 23266
rect 15036 22428 15316 22484
rect 15260 22370 15316 22428
rect 15260 22318 15262 22370
rect 15314 22318 15316 22370
rect 15260 22306 15316 22318
rect 16044 22372 16100 22382
rect 15932 22258 15988 22270
rect 15932 22206 15934 22258
rect 15986 22206 15988 22258
rect 15036 22148 15092 22158
rect 14924 22146 15092 22148
rect 14924 22094 15038 22146
rect 15090 22094 15092 22146
rect 14924 22092 15092 22094
rect 15036 22082 15092 22092
rect 15518 21980 15782 21990
rect 15574 21924 15622 21980
rect 15678 21924 15726 21980
rect 15518 21914 15782 21924
rect 15932 21476 15988 22206
rect 16044 21586 16100 22316
rect 16044 21534 16046 21586
rect 16098 21534 16100 21586
rect 16044 21522 16100 21534
rect 14588 20638 14590 20690
rect 14642 20638 14644 20690
rect 14588 20626 14644 20638
rect 15260 20804 15316 20814
rect 15036 20580 15092 20590
rect 15036 20578 15204 20580
rect 15036 20526 15038 20578
rect 15090 20526 15204 20578
rect 15036 20524 15204 20526
rect 15036 20514 15092 20524
rect 15148 20132 15204 20524
rect 15148 20066 15204 20076
rect 14812 20018 14868 20030
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14140 18610 14196 18620
rect 14252 19234 14308 19246
rect 14252 19182 14254 19234
rect 14306 19182 14308 19234
rect 14028 17666 14084 17678
rect 14028 17614 14030 17666
rect 14082 17614 14084 17666
rect 13916 15876 13972 15886
rect 13916 15314 13972 15820
rect 13916 15262 13918 15314
rect 13970 15262 13972 15314
rect 13916 15250 13972 15262
rect 14028 15316 14084 17614
rect 14140 15316 14196 15326
rect 14028 15260 14140 15316
rect 14140 15222 14196 15260
rect 14252 15202 14308 19182
rect 14364 19124 14420 19134
rect 14364 17220 14420 19068
rect 14812 18674 14868 19966
rect 15036 19460 15092 19470
rect 15148 19460 15204 19470
rect 15036 19458 15148 19460
rect 15036 19406 15038 19458
rect 15090 19406 15148 19458
rect 15036 19404 15148 19406
rect 15036 19394 15092 19404
rect 14812 18622 14814 18674
rect 14866 18622 14868 18674
rect 14812 18610 14868 18622
rect 14700 18564 14756 18574
rect 14700 18470 14756 18508
rect 15036 17892 15092 17902
rect 15036 17778 15092 17836
rect 15036 17726 15038 17778
rect 15090 17726 15092 17778
rect 15036 17714 15092 17726
rect 15148 17666 15204 19404
rect 15260 18788 15316 20748
rect 15518 20412 15782 20422
rect 15574 20356 15622 20412
rect 15678 20356 15726 20412
rect 15518 20346 15782 20356
rect 15484 20132 15540 20142
rect 15484 19684 15540 20076
rect 15820 20132 15876 20142
rect 15484 19618 15540 19628
rect 15596 20020 15652 20030
rect 15596 19346 15652 19964
rect 15820 19908 15876 20076
rect 15932 20020 15988 21420
rect 16044 21364 16100 21374
rect 16044 21270 16100 21308
rect 16044 20802 16100 20814
rect 16044 20750 16046 20802
rect 16098 20750 16100 20802
rect 16044 20692 16100 20750
rect 16044 20626 16100 20636
rect 15932 19964 16100 20020
rect 15820 19906 15988 19908
rect 15820 19854 15822 19906
rect 15874 19854 15988 19906
rect 15820 19852 15988 19854
rect 15820 19842 15876 19852
rect 15596 19294 15598 19346
rect 15650 19294 15652 19346
rect 15596 19282 15652 19294
rect 15708 19236 15764 19246
rect 15708 19142 15764 19180
rect 15518 18844 15782 18854
rect 15574 18788 15622 18844
rect 15678 18788 15726 18844
rect 15518 18778 15782 18788
rect 15260 18722 15316 18732
rect 15484 18676 15540 18686
rect 15372 18620 15484 18676
rect 15148 17614 15150 17666
rect 15202 17614 15204 17666
rect 15148 17602 15204 17614
rect 15260 18564 15316 18574
rect 15260 17444 15316 18508
rect 14364 17154 14420 17164
rect 15148 17388 15316 17444
rect 14588 17108 14644 17118
rect 14588 16882 14644 17052
rect 14588 16830 14590 16882
rect 14642 16830 14644 16882
rect 14588 16818 14644 16830
rect 15036 16882 15092 16894
rect 15036 16830 15038 16882
rect 15090 16830 15092 16882
rect 14476 15988 14532 15998
rect 14476 15894 14532 15932
rect 15036 15876 15092 16830
rect 15036 15782 15092 15820
rect 15148 15652 15204 17388
rect 15036 15596 15204 15652
rect 15260 16098 15316 16110
rect 15260 16046 15262 16098
rect 15314 16046 15316 16098
rect 14252 15150 14254 15202
rect 14306 15150 14308 15202
rect 13804 15092 14196 15148
rect 14252 15138 14308 15150
rect 14924 15316 14980 15326
rect 13580 14590 13582 14642
rect 13634 14590 13636 14642
rect 13580 14578 13636 14590
rect 13804 14644 13860 14654
rect 13804 13970 13860 14588
rect 13804 13918 13806 13970
rect 13858 13918 13860 13970
rect 13804 13906 13860 13918
rect 13580 12738 13636 12750
rect 13580 12686 13582 12738
rect 13634 12686 13636 12738
rect 13580 12404 13636 12686
rect 13580 12338 13636 12348
rect 14140 12402 14196 15092
rect 14252 14868 14308 14878
rect 14308 14812 14420 14868
rect 14252 14802 14308 14812
rect 14252 14420 14308 14430
rect 14252 14326 14308 14364
rect 14364 14420 14420 14812
rect 14588 14420 14644 14430
rect 14364 14418 14644 14420
rect 14364 14366 14590 14418
rect 14642 14366 14644 14418
rect 14364 14364 14644 14366
rect 14252 13076 14308 13086
rect 14364 13076 14420 14364
rect 14588 14354 14644 14364
rect 14700 13858 14756 13870
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13300 14756 13806
rect 14700 13234 14756 13244
rect 14252 13074 14420 13076
rect 14252 13022 14254 13074
rect 14306 13022 14420 13074
rect 14252 13020 14420 13022
rect 14252 13010 14308 13020
rect 14140 12350 14142 12402
rect 14194 12350 14196 12402
rect 14140 12338 14196 12350
rect 14364 12404 14420 13020
rect 14812 12964 14868 12974
rect 14364 12338 14420 12348
rect 14588 12962 14868 12964
rect 14588 12910 14814 12962
rect 14866 12910 14868 12962
rect 14588 12908 14868 12910
rect 13692 12068 13748 12078
rect 13692 12066 13860 12068
rect 13692 12014 13694 12066
rect 13746 12014 13860 12066
rect 13692 12012 13860 12014
rect 13692 12002 13748 12012
rect 13692 11508 13748 11518
rect 13692 11414 13748 11452
rect 13580 11172 13636 11182
rect 13468 10722 13524 10734
rect 13468 10670 13470 10722
rect 13522 10670 13524 10722
rect 13356 10612 13412 10622
rect 13468 10612 13524 10670
rect 13580 10722 13636 11116
rect 13580 10670 13582 10722
rect 13634 10670 13636 10722
rect 13580 10658 13636 10670
rect 13412 10556 13524 10612
rect 13356 10546 13412 10556
rect 13804 10498 13860 12012
rect 14476 11954 14532 11966
rect 14476 11902 14478 11954
rect 14530 11902 14532 11954
rect 14140 11508 14196 11518
rect 14140 11414 14196 11452
rect 14476 11396 14532 11902
rect 14588 11844 14644 12908
rect 14812 12898 14868 12908
rect 14924 12178 14980 15260
rect 15036 13860 15092 15596
rect 15036 13766 15092 13804
rect 15148 15428 15204 15438
rect 14924 12126 14926 12178
rect 14978 12126 14980 12178
rect 14924 12114 14980 12126
rect 15036 13300 15092 13310
rect 15036 12290 15092 13244
rect 15036 12238 15038 12290
rect 15090 12238 15092 12290
rect 14588 11506 14644 11788
rect 14588 11454 14590 11506
rect 14642 11454 14644 11506
rect 14588 11442 14644 11454
rect 14812 11956 14868 11966
rect 14252 11340 14532 11396
rect 14140 11172 14196 11182
rect 14252 11172 14308 11340
rect 14196 11116 14308 11172
rect 14364 11172 14420 11182
rect 14140 10722 14196 11116
rect 14140 10670 14142 10722
rect 14194 10670 14196 10722
rect 14140 10658 14196 10670
rect 13804 10446 13806 10498
rect 13858 10446 13860 10498
rect 13692 9940 13748 9950
rect 13356 8930 13412 8942
rect 13356 8878 13358 8930
rect 13410 8878 13412 8930
rect 13356 8820 13412 8878
rect 13412 8764 13524 8820
rect 13356 8754 13412 8764
rect 13468 8258 13524 8764
rect 13468 8206 13470 8258
rect 13522 8206 13524 8258
rect 13468 8194 13524 8206
rect 13580 8260 13636 8270
rect 13692 8260 13748 9884
rect 13804 9828 13860 10446
rect 14364 10610 14420 11116
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14364 10500 14420 10558
rect 14588 10610 14644 10622
rect 14588 10558 14590 10610
rect 14642 10558 14644 10610
rect 14364 10434 14420 10444
rect 14476 10498 14532 10510
rect 14476 10446 14478 10498
rect 14530 10446 14532 10498
rect 14476 10276 14532 10446
rect 13916 10220 14532 10276
rect 14588 10388 14644 10558
rect 14700 10612 14756 10622
rect 14700 10518 14756 10556
rect 13916 10050 13972 10220
rect 13916 9998 13918 10050
rect 13970 9998 13972 10050
rect 13916 9986 13972 9998
rect 14252 9940 14308 9950
rect 14588 9940 14644 10332
rect 14252 9846 14308 9884
rect 14476 9884 14644 9940
rect 13804 9156 13860 9772
rect 14476 9828 14532 9884
rect 14476 9604 14532 9772
rect 14700 9604 14756 9614
rect 14476 9602 14756 9604
rect 14476 9550 14702 9602
rect 14754 9550 14756 9602
rect 14476 9548 14756 9550
rect 14700 9538 14756 9548
rect 13804 9062 13860 9100
rect 14700 9380 14756 9390
rect 14700 9154 14756 9324
rect 14700 9102 14702 9154
rect 14754 9102 14756 9154
rect 14700 9090 14756 9102
rect 14476 9042 14532 9054
rect 14476 8990 14478 9042
rect 14530 8990 14532 9042
rect 14476 8820 14532 8990
rect 14476 8754 14532 8764
rect 13916 8260 13972 8270
rect 13692 8258 13972 8260
rect 13692 8206 13918 8258
rect 13970 8206 13972 8258
rect 13692 8204 13972 8206
rect 13580 8036 13636 8204
rect 13692 8036 13748 8046
rect 13580 8034 13748 8036
rect 13580 7982 13694 8034
rect 13746 7982 13748 8034
rect 13580 7980 13748 7982
rect 13692 7970 13748 7980
rect 13804 8034 13860 8046
rect 13804 7982 13806 8034
rect 13858 7982 13860 8034
rect 13132 7858 13188 7868
rect 12908 7700 12964 7710
rect 12124 7588 12180 7598
rect 12124 7494 12180 7532
rect 11228 7476 11284 7486
rect 11228 7382 11284 7420
rect 11900 7476 11956 7486
rect 12572 7476 12628 7486
rect 11900 7382 11956 7420
rect 12236 7474 12628 7476
rect 12236 7422 12574 7474
rect 12626 7422 12628 7474
rect 12236 7420 12628 7422
rect 12236 7362 12292 7420
rect 12572 7410 12628 7420
rect 12908 7474 12964 7644
rect 13804 7700 13860 7982
rect 13804 7634 13860 7644
rect 13916 7588 13972 8204
rect 14140 8146 14196 8158
rect 14140 8094 14142 8146
rect 14194 8094 14196 8146
rect 14028 7588 14084 7598
rect 13972 7586 14084 7588
rect 13972 7534 14030 7586
rect 14082 7534 14084 7586
rect 13972 7532 14084 7534
rect 13916 7494 13972 7532
rect 14028 7522 14084 7532
rect 12908 7422 12910 7474
rect 12962 7422 12964 7474
rect 12908 7410 12964 7422
rect 14140 7476 14196 8094
rect 14588 7476 14644 7486
rect 14196 7474 14644 7476
rect 14196 7422 14590 7474
rect 14642 7422 14644 7474
rect 14196 7420 14644 7422
rect 14140 7382 14196 7420
rect 12236 7310 12238 7362
rect 12290 7310 12292 7362
rect 12236 7298 12292 7310
rect 13356 7362 13412 7374
rect 13356 7310 13358 7362
rect 13410 7310 13412 7362
rect 9996 6066 10052 6076
rect 10444 6076 11060 6132
rect 8204 5906 8260 5918
rect 8204 5854 8206 5906
rect 8258 5854 8260 5906
rect 8092 5236 8148 5246
rect 8092 5122 8148 5180
rect 8204 5234 8260 5854
rect 8316 5908 8372 5918
rect 8316 5814 8372 5852
rect 8764 5908 8820 5918
rect 8764 5814 8820 5852
rect 10220 5906 10276 5918
rect 10220 5854 10222 5906
rect 10274 5854 10276 5906
rect 10108 5796 10164 5806
rect 8365 5516 8629 5526
rect 8421 5460 8469 5516
rect 8525 5460 8573 5516
rect 8365 5450 8629 5460
rect 8204 5182 8206 5234
rect 8258 5182 8260 5234
rect 8204 5170 8260 5182
rect 8092 5070 8094 5122
rect 8146 5070 8148 5122
rect 8092 5058 8148 5070
rect 8316 5124 8372 5134
rect 8316 5030 8372 5068
rect 8764 5124 8820 5134
rect 9212 5124 9268 5134
rect 8764 5122 9492 5124
rect 8764 5070 8766 5122
rect 8818 5070 9214 5122
rect 9266 5070 9492 5122
rect 8764 5068 9492 5070
rect 8764 5058 8820 5068
rect 9212 5058 9268 5068
rect 9436 4564 9492 5068
rect 9548 5012 9604 5022
rect 9548 4918 9604 4956
rect 9548 4564 9604 4574
rect 9436 4562 9604 4564
rect 9436 4510 9550 4562
rect 9602 4510 9604 4562
rect 9436 4508 9604 4510
rect 9548 4498 9604 4508
rect 9772 4564 9828 4574
rect 9772 4470 9828 4508
rect 8204 4452 8260 4462
rect 8204 4358 8260 4396
rect 9884 4452 9940 4462
rect 10108 4452 10164 5740
rect 10220 5236 10276 5854
rect 10444 5906 10500 6076
rect 10444 5854 10446 5906
rect 10498 5854 10500 5906
rect 10444 5842 10500 5854
rect 10668 5906 10724 5918
rect 10668 5854 10670 5906
rect 10722 5854 10724 5906
rect 10556 5794 10612 5806
rect 10556 5742 10558 5794
rect 10610 5742 10612 5794
rect 10556 5236 10612 5742
rect 10668 5796 10724 5854
rect 10668 5730 10724 5740
rect 10780 5236 10836 5246
rect 10556 5180 10724 5236
rect 10220 5170 10276 5180
rect 9884 4450 10612 4452
rect 9884 4398 9886 4450
rect 9938 4398 10612 4450
rect 9884 4396 10612 4398
rect 9884 4386 9940 4396
rect 7980 4286 7982 4338
rect 8034 4286 8036 4338
rect 7980 4274 8036 4286
rect 10556 4338 10612 4396
rect 10556 4286 10558 4338
rect 10610 4286 10612 4338
rect 10556 4274 10612 4286
rect 10668 4340 10724 5180
rect 10780 5142 10836 5180
rect 10892 5124 10948 5134
rect 10892 5030 10948 5068
rect 10668 4274 10724 4284
rect 11004 4564 11060 6076
rect 12684 5908 12740 5918
rect 11676 5348 11732 5358
rect 11676 5254 11732 5292
rect 12684 5348 12740 5852
rect 11004 4338 11060 4508
rect 11788 5236 11844 5246
rect 11788 4452 11844 5180
rect 12684 5234 12740 5292
rect 12684 5182 12686 5234
rect 12738 5182 12740 5234
rect 12684 5170 12740 5182
rect 13356 5236 13412 7310
rect 14588 7140 14644 7420
rect 14588 7074 14644 7084
rect 14812 6020 14868 11900
rect 14924 11844 14980 11854
rect 14924 8820 14980 11788
rect 15036 10612 15092 12238
rect 15148 10724 15204 15372
rect 15260 14532 15316 16046
rect 15260 14466 15316 14476
rect 15372 13748 15428 18620
rect 15484 18610 15540 18620
rect 15820 18452 15876 18462
rect 15932 18452 15988 19852
rect 16044 19236 16100 19964
rect 16156 19460 16212 23214
rect 16268 22372 16324 23884
rect 16268 22306 16324 22316
rect 16492 23154 16548 23166
rect 16492 23102 16494 23154
rect 16546 23102 16548 23154
rect 16268 22148 16324 22158
rect 16268 21586 16324 22092
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 16268 21522 16324 21534
rect 16268 21364 16324 21374
rect 16268 20130 16324 21308
rect 16268 20078 16270 20130
rect 16322 20078 16324 20130
rect 16268 20066 16324 20078
rect 16492 20132 16548 23102
rect 16604 22148 16660 25230
rect 16828 24388 16884 24398
rect 16604 22082 16660 22092
rect 16716 23938 16772 23950
rect 16716 23886 16718 23938
rect 16770 23886 16772 23938
rect 16716 23380 16772 23886
rect 16604 21812 16660 21822
rect 16604 20690 16660 21756
rect 16604 20638 16606 20690
rect 16658 20638 16660 20690
rect 16604 20468 16660 20638
rect 16716 20692 16772 23324
rect 16716 20626 16772 20636
rect 16716 20468 16772 20478
rect 16604 20412 16716 20468
rect 16716 20402 16772 20412
rect 16828 20242 16884 24332
rect 17276 23940 17332 23950
rect 16940 23380 16996 23390
rect 16940 23286 16996 23324
rect 16940 22596 16996 22606
rect 16940 21364 16996 22540
rect 17276 22370 17332 23884
rect 17388 23380 17444 25452
rect 17500 24722 17556 26236
rect 19180 26290 19236 26302
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 19068 26066 19124 26078
rect 19068 26014 19070 26066
rect 19122 26014 19124 26066
rect 17612 25508 17668 25518
rect 17612 25414 17668 25452
rect 19068 25508 19124 26014
rect 19180 26068 19236 26238
rect 19628 26180 19684 26190
rect 19628 26086 19684 26124
rect 20076 26178 20132 26190
rect 20076 26126 20078 26178
rect 20130 26126 20132 26178
rect 19180 26002 19236 26012
rect 19964 26068 20020 26078
rect 18732 25396 18788 25406
rect 17500 24670 17502 24722
rect 17554 24670 17556 24722
rect 17500 24658 17556 24670
rect 18060 25284 18116 25294
rect 17500 24500 17556 24510
rect 17500 24406 17556 24444
rect 17948 23940 18004 23950
rect 17388 23324 17780 23380
rect 17612 23044 17668 23054
rect 17276 22318 17278 22370
rect 17330 22318 17332 22370
rect 17276 22306 17332 22318
rect 17500 23042 17668 23044
rect 17500 22990 17614 23042
rect 17666 22990 17668 23042
rect 17500 22988 17668 22990
rect 16940 21298 16996 21308
rect 17052 20804 17108 20814
rect 17052 20710 17108 20748
rect 16828 20190 16830 20242
rect 16882 20190 16884 20242
rect 16828 20178 16884 20190
rect 16716 20132 16772 20142
rect 16492 20066 16548 20076
rect 16604 20076 16716 20132
rect 16492 19908 16548 19918
rect 16604 19908 16660 20076
rect 16716 20066 16772 20076
rect 17388 20020 17444 20030
rect 16492 19906 16660 19908
rect 16492 19854 16494 19906
rect 16546 19854 16660 19906
rect 16492 19852 16660 19854
rect 16492 19842 16548 19852
rect 16156 19394 16212 19404
rect 16492 19572 16548 19582
rect 16044 19180 16324 19236
rect 15820 18450 15988 18452
rect 15820 18398 15822 18450
rect 15874 18398 15988 18450
rect 15820 18396 15988 18398
rect 15820 18386 15876 18396
rect 15820 18228 15876 18238
rect 15820 17554 15876 18172
rect 16156 18228 16212 18238
rect 16156 18134 16212 18172
rect 15820 17502 15822 17554
rect 15874 17502 15876 17554
rect 15820 17490 15876 17502
rect 15518 17276 15782 17286
rect 15574 17220 15622 17276
rect 15678 17220 15726 17276
rect 15518 17210 15782 17220
rect 15596 16996 15652 17006
rect 16268 16996 16324 19180
rect 16492 19122 16548 19516
rect 16492 19070 16494 19122
rect 16546 19070 16548 19122
rect 16492 18564 16548 19070
rect 16604 18676 16660 19852
rect 17052 20018 17444 20020
rect 17052 19966 17390 20018
rect 17442 19966 17444 20018
rect 17052 19964 17444 19966
rect 16604 18610 16660 18620
rect 16940 19346 16996 19358
rect 16940 19294 16942 19346
rect 16994 19294 16996 19346
rect 16492 18498 16548 18508
rect 15596 16902 15652 16940
rect 16156 16940 16324 16996
rect 16828 18452 16884 18462
rect 15518 15708 15782 15718
rect 15574 15652 15622 15708
rect 15678 15652 15726 15708
rect 15518 15642 15782 15652
rect 15484 15428 15540 15438
rect 15484 15334 15540 15372
rect 16044 15428 16100 15438
rect 16156 15428 16212 16940
rect 16604 16660 16660 16670
rect 16604 16566 16660 16604
rect 16604 15986 16660 15998
rect 16604 15934 16606 15986
rect 16658 15934 16660 15986
rect 16268 15876 16324 15886
rect 16268 15874 16436 15876
rect 16268 15822 16270 15874
rect 16322 15822 16436 15874
rect 16268 15820 16436 15822
rect 16268 15810 16324 15820
rect 16044 15426 16212 15428
rect 16044 15374 16046 15426
rect 16098 15374 16212 15426
rect 16044 15372 16212 15374
rect 16268 15428 16324 15438
rect 16044 15362 16100 15372
rect 16268 15314 16324 15372
rect 16268 15262 16270 15314
rect 16322 15262 16324 15314
rect 16268 15250 16324 15262
rect 16380 15316 16436 15820
rect 16380 15222 16436 15260
rect 16492 15874 16548 15886
rect 16492 15822 16494 15874
rect 16546 15822 16548 15874
rect 16156 15204 16212 15214
rect 16156 15092 16324 15148
rect 16044 14532 16100 14542
rect 16100 14476 16212 14532
rect 16044 14438 16100 14476
rect 16044 14308 16100 14318
rect 15518 14140 15782 14150
rect 15574 14084 15622 14140
rect 15678 14084 15726 14140
rect 15518 14074 15782 14084
rect 15708 13972 15764 13982
rect 15708 13878 15764 13916
rect 15596 13860 15652 13870
rect 15372 13692 15540 13748
rect 15372 13524 15428 13534
rect 15372 13430 15428 13468
rect 15372 13076 15428 13086
rect 15484 13076 15540 13692
rect 15372 13074 15540 13076
rect 15372 13022 15374 13074
rect 15426 13022 15540 13074
rect 15372 13020 15540 13022
rect 15372 13010 15428 13020
rect 15484 12852 15540 12862
rect 15596 12852 15652 13804
rect 16044 13412 16100 14252
rect 16156 13746 16212 14476
rect 16268 14420 16324 15092
rect 16380 14420 16436 14430
rect 16268 14418 16436 14420
rect 16268 14366 16382 14418
rect 16434 14366 16436 14418
rect 16268 14364 16436 14366
rect 16156 13694 16158 13746
rect 16210 13694 16212 13746
rect 16156 13682 16212 13694
rect 16380 13748 16436 14364
rect 16492 13972 16548 15822
rect 16604 14420 16660 15934
rect 16828 15148 16884 18396
rect 16604 14084 16660 14364
rect 16716 15092 16884 15148
rect 16940 18340 16996 19294
rect 17052 19236 17108 19964
rect 17388 19954 17444 19964
rect 17500 20020 17556 22988
rect 17612 22978 17668 22988
rect 17724 21810 17780 23324
rect 17836 23044 17892 23054
rect 17836 22950 17892 22988
rect 17836 22596 17892 22606
rect 17836 22370 17892 22540
rect 17836 22318 17838 22370
rect 17890 22318 17892 22370
rect 17836 22306 17892 22318
rect 17724 21758 17726 21810
rect 17778 21758 17780 21810
rect 17724 21746 17780 21758
rect 17612 21586 17668 21598
rect 17612 21534 17614 21586
rect 17666 21534 17668 21586
rect 17612 21476 17668 21534
rect 17948 21586 18004 23884
rect 18060 23268 18116 25228
rect 18396 24724 18452 24734
rect 18284 24610 18340 24622
rect 18284 24558 18286 24610
rect 18338 24558 18340 24610
rect 18060 23202 18116 23212
rect 18172 23826 18228 23838
rect 18172 23774 18174 23826
rect 18226 23774 18228 23826
rect 18172 22372 18228 23774
rect 18284 23380 18340 24558
rect 18396 23604 18452 24668
rect 18508 24276 18564 24286
rect 18508 23938 18564 24220
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18508 23874 18564 23886
rect 18396 23538 18452 23548
rect 18284 23324 18452 23380
rect 18284 23154 18340 23166
rect 18284 23102 18286 23154
rect 18338 23102 18340 23154
rect 18284 23044 18340 23102
rect 18284 22978 18340 22988
rect 18172 22316 18340 22372
rect 17948 21534 17950 21586
rect 18002 21534 18004 21586
rect 17948 21522 18004 21534
rect 18172 22148 18228 22158
rect 17612 21410 17668 21420
rect 17612 20020 17668 20030
rect 17500 19964 17612 20020
rect 17052 19142 17108 19180
rect 17276 19684 17332 19694
rect 16716 14308 16772 15092
rect 16940 14868 16996 18284
rect 17276 17780 17332 19628
rect 17500 19460 17556 19964
rect 17612 19954 17668 19964
rect 17500 19394 17556 19404
rect 17612 19234 17668 19246
rect 17612 19182 17614 19234
rect 17666 19182 17668 19234
rect 17388 18452 17444 18462
rect 17388 18358 17444 18396
rect 17388 17780 17444 17790
rect 17276 17778 17444 17780
rect 17276 17726 17390 17778
rect 17442 17726 17444 17778
rect 17276 17724 17444 17726
rect 17388 16882 17444 17724
rect 17500 17780 17556 17790
rect 17612 17780 17668 19182
rect 18172 19122 18228 22092
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 19058 18228 19070
rect 18284 18564 18340 22316
rect 18396 22036 18452 23324
rect 18620 22932 18676 22942
rect 18620 22370 18676 22876
rect 18620 22318 18622 22370
rect 18674 22318 18676 22370
rect 18620 22306 18676 22318
rect 18396 21970 18452 21980
rect 18284 18498 18340 18508
rect 18508 20914 18564 20926
rect 18508 20862 18510 20914
rect 18562 20862 18564 20914
rect 18508 18900 18564 20862
rect 18396 18452 18452 18462
rect 18508 18452 18564 18844
rect 18396 18450 18564 18452
rect 18396 18398 18398 18450
rect 18450 18398 18564 18450
rect 18396 18396 18564 18398
rect 17724 18340 17780 18350
rect 18060 18340 18116 18350
rect 17780 18338 18116 18340
rect 17780 18286 18062 18338
rect 18114 18286 18116 18338
rect 17780 18284 18116 18286
rect 17724 18274 17780 18284
rect 18060 18274 18116 18284
rect 17612 17724 17780 17780
rect 17500 17668 17556 17724
rect 17500 17666 17668 17668
rect 17500 17614 17502 17666
rect 17554 17614 17668 17666
rect 17500 17612 17668 17614
rect 17500 17602 17556 17612
rect 17388 16830 17390 16882
rect 17442 16830 17444 16882
rect 17388 16818 17444 16830
rect 17612 16882 17668 17612
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 17612 16818 17668 16830
rect 16940 14802 16996 14812
rect 17164 16660 17220 16670
rect 17164 15986 17220 16604
rect 17724 16210 17780 17724
rect 18172 17668 18228 17678
rect 18172 17574 18228 17612
rect 18396 17444 18452 18396
rect 18396 17378 18452 17388
rect 18732 18340 18788 25340
rect 19068 24722 19124 25452
rect 19068 24670 19070 24722
rect 19122 24670 19124 24722
rect 19068 24658 19124 24670
rect 19740 25506 19796 25518
rect 19740 25454 19742 25506
rect 19794 25454 19796 25506
rect 19740 25396 19796 25454
rect 19740 23042 19796 25340
rect 19964 25396 20020 26012
rect 20076 25844 20132 26126
rect 21084 26180 21140 26190
rect 20076 25778 20132 25788
rect 20972 26066 21028 26078
rect 20972 26014 20974 26066
rect 21026 26014 21028 26066
rect 20188 25396 20244 25406
rect 19964 25394 20244 25396
rect 19964 25342 20190 25394
rect 20242 25342 20244 25394
rect 19964 25340 20244 25342
rect 19964 23940 20020 25340
rect 20188 25330 20244 25340
rect 20972 25396 21028 26014
rect 20972 25330 21028 25340
rect 20636 25282 20692 25294
rect 20636 25230 20638 25282
rect 20690 25230 20692 25282
rect 20412 24722 20468 24734
rect 20412 24670 20414 24722
rect 20466 24670 20468 24722
rect 20412 24388 20468 24670
rect 20412 24322 20468 24332
rect 20636 24724 20692 25230
rect 19964 23846 20020 23884
rect 20076 24052 20132 24062
rect 20636 24052 20692 24668
rect 20076 23380 20132 23996
rect 20412 23996 20692 24052
rect 19740 22990 19742 23042
rect 19794 22990 19796 23042
rect 19740 22978 19796 22990
rect 19852 23324 20132 23380
rect 20188 23380 20244 23390
rect 19628 22708 19684 22718
rect 19628 21698 19684 22652
rect 19628 21646 19630 21698
rect 19682 21646 19684 21698
rect 19628 21634 19684 21646
rect 19852 21586 19908 23324
rect 19852 21534 19854 21586
rect 19906 21534 19908 21586
rect 19852 21522 19908 21534
rect 19964 23154 20020 23166
rect 19964 23102 19966 23154
rect 20018 23102 20020 23154
rect 19404 19908 19460 19918
rect 19404 19346 19460 19852
rect 19404 19294 19406 19346
rect 19458 19294 19460 19346
rect 19404 19282 19460 19294
rect 19516 19906 19572 19918
rect 19516 19854 19518 19906
rect 19570 19854 19572 19906
rect 18844 18562 18900 18574
rect 18844 18510 18846 18562
rect 18898 18510 18900 18562
rect 18844 18452 18900 18510
rect 18844 18386 18900 18396
rect 19292 18564 19348 18574
rect 18732 16884 18788 18284
rect 19292 17668 19348 18508
rect 19516 18116 19572 19854
rect 19628 19012 19684 19022
rect 19628 18918 19684 18956
rect 19740 18900 19796 18910
rect 19740 18788 19796 18844
rect 18732 16818 18788 16828
rect 18844 17666 19348 17668
rect 18844 17614 19294 17666
rect 19346 17614 19348 17666
rect 18844 17612 19348 17614
rect 17724 16158 17726 16210
rect 17778 16158 17780 16210
rect 17724 16146 17780 16158
rect 17164 15934 17166 15986
rect 17218 15934 17220 15986
rect 17164 14420 17220 15934
rect 17948 16098 18004 16110
rect 18732 16100 18788 16110
rect 17948 16046 17950 16098
rect 18002 16046 18004 16098
rect 17724 15314 17780 15326
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 17724 15204 17780 15262
rect 17724 15138 17780 15148
rect 17164 14326 17220 14364
rect 16716 14242 16772 14252
rect 16604 14018 16660 14028
rect 16940 14084 16996 14094
rect 16492 13906 16548 13916
rect 16716 13860 16772 13898
rect 16716 13794 16772 13804
rect 16380 13692 16660 13748
rect 15484 12850 15652 12852
rect 15484 12798 15486 12850
rect 15538 12798 15652 12850
rect 15484 12796 15652 12798
rect 15932 13356 16100 13412
rect 16492 13524 16548 13534
rect 15932 12850 15988 13356
rect 16268 13076 16324 13086
rect 16492 13076 16548 13468
rect 16268 13074 16548 13076
rect 16268 13022 16270 13074
rect 16322 13022 16548 13074
rect 16268 13020 16548 13022
rect 16268 13010 16324 13020
rect 16604 12964 16660 13692
rect 15932 12798 15934 12850
rect 15986 12798 15988 12850
rect 15484 12786 15540 12796
rect 15260 12738 15316 12750
rect 15260 12686 15262 12738
rect 15314 12686 15316 12738
rect 15260 11508 15316 12686
rect 15518 12572 15782 12582
rect 15574 12516 15622 12572
rect 15678 12516 15726 12572
rect 15518 12506 15782 12516
rect 15820 12404 15876 12414
rect 15932 12404 15988 12798
rect 16380 12908 16604 12964
rect 16380 12850 16436 12908
rect 16604 12898 16660 12908
rect 16380 12798 16382 12850
rect 16434 12798 16436 12850
rect 16380 12786 16436 12798
rect 15820 12402 15988 12404
rect 15820 12350 15822 12402
rect 15874 12350 15988 12402
rect 15820 12348 15988 12350
rect 16156 12738 16212 12750
rect 16156 12686 16158 12738
rect 16210 12686 16212 12738
rect 15820 12338 15876 12348
rect 15260 11442 15316 11452
rect 15372 11620 15428 11630
rect 15260 11284 15316 11294
rect 15372 11284 15428 11564
rect 16156 11620 16212 12686
rect 16380 12404 16436 12414
rect 16380 12310 16436 12348
rect 16940 11956 16996 14028
rect 17388 13972 17444 13982
rect 17388 13878 17444 13916
rect 17612 13860 17668 13870
rect 17612 13746 17668 13804
rect 17612 13694 17614 13746
rect 17666 13694 17668 13746
rect 17612 13682 17668 13694
rect 17948 13748 18004 16046
rect 18508 16098 18788 16100
rect 18508 16046 18734 16098
rect 18786 16046 18788 16098
rect 18508 16044 18788 16046
rect 18060 15988 18116 15998
rect 18060 15426 18116 15932
rect 18060 15374 18062 15426
rect 18114 15374 18116 15426
rect 18060 15148 18116 15374
rect 18508 15148 18564 16044
rect 18732 16034 18788 16044
rect 18844 16100 18900 17612
rect 19292 17602 19348 17612
rect 19404 18060 19572 18116
rect 19628 18732 19796 18788
rect 19404 17332 19460 18060
rect 19292 16884 19348 16894
rect 19292 16790 19348 16828
rect 18844 15876 18900 16044
rect 18620 15820 18900 15876
rect 18620 15314 18676 15820
rect 18620 15262 18622 15314
rect 18674 15262 18676 15314
rect 18620 15250 18676 15262
rect 18732 15538 18788 15550
rect 18732 15486 18734 15538
rect 18786 15486 18788 15538
rect 18732 15316 18788 15486
rect 19180 15316 19236 15326
rect 18732 15314 19236 15316
rect 18732 15262 19182 15314
rect 19234 15262 19236 15314
rect 18732 15260 19236 15262
rect 19180 15250 19236 15260
rect 18060 15092 18452 15148
rect 18508 15092 18788 15148
rect 18172 14868 18228 14878
rect 18228 14812 18340 14868
rect 18172 14802 18228 14812
rect 18172 14532 18228 14542
rect 17948 13186 18004 13692
rect 17948 13134 17950 13186
rect 18002 13134 18004 13186
rect 17948 13122 18004 13134
rect 18060 14530 18228 14532
rect 18060 14478 18174 14530
rect 18226 14478 18228 14530
rect 18060 14476 18228 14478
rect 16940 11890 16996 11900
rect 17052 13076 17108 13086
rect 17052 12850 17108 13020
rect 17052 12798 17054 12850
rect 17106 12798 17108 12850
rect 16156 11554 16212 11564
rect 15260 11282 15428 11284
rect 15260 11230 15262 11282
rect 15314 11230 15428 11282
rect 15260 11228 15428 11230
rect 15260 10948 15316 11228
rect 15708 11172 15764 11182
rect 15260 10882 15316 10892
rect 15372 11170 15764 11172
rect 15372 11118 15710 11170
rect 15762 11118 15764 11170
rect 15372 11116 15764 11118
rect 15372 10836 15428 11116
rect 15708 11106 15764 11116
rect 15518 11004 15782 11014
rect 15574 10948 15622 11004
rect 15678 10948 15726 11004
rect 15518 10938 15782 10948
rect 15484 10836 15540 10846
rect 15372 10834 15540 10836
rect 15372 10782 15486 10834
rect 15538 10782 15540 10834
rect 15372 10780 15540 10782
rect 15148 10658 15204 10668
rect 15036 10388 15092 10556
rect 15372 10610 15428 10622
rect 15372 10558 15374 10610
rect 15426 10558 15428 10610
rect 15372 10500 15428 10558
rect 15484 10612 15540 10780
rect 16604 10724 16660 10734
rect 16604 10630 16660 10668
rect 15484 10546 15540 10556
rect 15708 10610 15764 10622
rect 15708 10558 15710 10610
rect 15762 10558 15764 10610
rect 15372 10434 15428 10444
rect 15708 10388 15764 10558
rect 16268 10612 16324 10622
rect 16044 10388 16100 10398
rect 15708 10332 16044 10388
rect 15036 10322 15092 10332
rect 16044 10294 16100 10332
rect 15372 9938 15428 9950
rect 15372 9886 15374 9938
rect 15426 9886 15428 9938
rect 15148 8932 15204 8942
rect 15372 8932 15428 9886
rect 15708 9828 15764 9838
rect 16156 9828 16212 9838
rect 15764 9772 15988 9828
rect 15708 9734 15764 9772
rect 15518 9436 15782 9446
rect 15574 9380 15622 9436
rect 15678 9380 15726 9436
rect 15518 9370 15782 9380
rect 15148 8930 15428 8932
rect 15148 8878 15150 8930
rect 15202 8878 15428 8930
rect 15148 8876 15428 8878
rect 15596 9156 15652 9166
rect 15148 8866 15204 8876
rect 14924 8370 14980 8764
rect 14924 8318 14926 8370
rect 14978 8318 14980 8370
rect 14924 8148 14980 8318
rect 14924 8082 14980 8092
rect 15260 8034 15316 8876
rect 15484 8596 15540 8606
rect 15484 8146 15540 8540
rect 15484 8094 15486 8146
rect 15538 8094 15540 8146
rect 15484 8082 15540 8094
rect 15596 8260 15652 9100
rect 15932 8596 15988 9772
rect 16156 9734 16212 9772
rect 16268 9604 16324 10556
rect 17052 10500 17108 12798
rect 17388 12964 17444 12974
rect 17612 12964 17668 12974
rect 17388 12850 17444 12908
rect 17388 12798 17390 12850
rect 17442 12798 17444 12850
rect 17388 12786 17444 12798
rect 17500 12962 17668 12964
rect 17500 12910 17614 12962
rect 17666 12910 17668 12962
rect 17500 12908 17668 12910
rect 17500 11172 17556 12908
rect 17612 12898 17668 12908
rect 18060 12292 18116 14476
rect 18172 14466 18228 14476
rect 18172 13972 18228 13982
rect 18284 13972 18340 14812
rect 18396 14644 18452 15092
rect 18620 14868 18676 14878
rect 18396 14588 18564 14644
rect 18172 13970 18284 13972
rect 18172 13918 18174 13970
rect 18226 13918 18284 13970
rect 18172 13916 18284 13918
rect 18172 13906 18228 13916
rect 18284 13878 18340 13916
rect 18396 14420 18452 14430
rect 18396 13860 18452 14364
rect 17724 12236 18116 12292
rect 18172 12852 18228 12862
rect 17612 12068 17668 12078
rect 17612 11974 17668 12012
rect 17500 11106 17556 11116
rect 17388 10724 17444 10734
rect 17388 10630 17444 10668
rect 17612 10612 17668 10622
rect 17724 10612 17780 12236
rect 18060 12068 18116 12078
rect 18172 12068 18228 12796
rect 18060 12066 18228 12068
rect 18060 12014 18062 12066
rect 18114 12014 18228 12066
rect 18060 12012 18228 12014
rect 18284 12292 18340 12302
rect 18060 11844 18116 12012
rect 18060 11778 18116 11788
rect 18284 10724 18340 12236
rect 18396 12290 18452 13804
rect 18508 13636 18564 14588
rect 18620 14530 18676 14812
rect 18732 14642 18788 15092
rect 18956 14868 19012 14878
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18732 14578 18788 14590
rect 18844 14812 18956 14868
rect 18620 14478 18622 14530
rect 18674 14478 18676 14530
rect 18620 14466 18676 14478
rect 18620 13636 18676 13646
rect 18508 13634 18676 13636
rect 18508 13582 18622 13634
rect 18674 13582 18676 13634
rect 18508 13580 18676 13582
rect 18508 12852 18564 13580
rect 18620 13570 18676 13580
rect 18732 13522 18788 13534
rect 18732 13470 18734 13522
rect 18786 13470 18788 13522
rect 18620 12964 18676 12974
rect 18620 12870 18676 12908
rect 18508 12758 18564 12796
rect 18508 12404 18564 12414
rect 18508 12310 18564 12348
rect 18732 12402 18788 13470
rect 18732 12350 18734 12402
rect 18786 12350 18788 12402
rect 18732 12338 18788 12350
rect 18844 12404 18900 14812
rect 18956 14802 19012 14812
rect 19404 14644 19460 17276
rect 19516 17890 19572 17902
rect 19516 17838 19518 17890
rect 19570 17838 19572 17890
rect 19516 16884 19572 17838
rect 19516 15314 19572 16828
rect 19516 15262 19518 15314
rect 19570 15262 19572 15314
rect 19516 15250 19572 15262
rect 19628 15148 19684 18732
rect 19740 18562 19796 18574
rect 19740 18510 19742 18562
rect 19794 18510 19796 18562
rect 19740 16772 19796 18510
rect 19964 17892 20020 23102
rect 20188 22482 20244 23324
rect 20188 22430 20190 22482
rect 20242 22430 20244 22482
rect 20188 22418 20244 22430
rect 20412 22370 20468 23996
rect 20412 22318 20414 22370
rect 20466 22318 20468 22370
rect 20412 22306 20468 22318
rect 20524 23826 20580 23838
rect 20524 23774 20526 23826
rect 20578 23774 20580 23826
rect 20412 21588 20468 21598
rect 20412 21494 20468 21532
rect 20412 20802 20468 20814
rect 20412 20750 20414 20802
rect 20466 20750 20468 20802
rect 20412 17892 20468 20750
rect 20524 20244 20580 23774
rect 20636 23828 20692 23838
rect 20636 23734 20692 23772
rect 20860 23714 20916 23726
rect 20860 23662 20862 23714
rect 20914 23662 20916 23714
rect 20860 22708 20916 23662
rect 21084 23042 21140 26124
rect 21532 25506 21588 26348
rect 22092 26404 22148 26414
rect 22092 26290 22148 26348
rect 26684 26402 26740 26460
rect 26684 26350 26686 26402
rect 26738 26350 26740 26402
rect 22092 26238 22094 26290
rect 22146 26238 22148 26290
rect 22092 26226 22148 26238
rect 22652 26292 22708 26302
rect 22652 26198 22708 26236
rect 21532 25454 21534 25506
rect 21586 25454 21588 25506
rect 21532 25442 21588 25454
rect 21980 26178 22036 26190
rect 21980 26126 21982 26178
rect 22034 26126 22036 26178
rect 21308 25396 21364 25406
rect 21308 25302 21364 25340
rect 21420 24834 21476 24846
rect 21420 24782 21422 24834
rect 21474 24782 21476 24834
rect 21196 24612 21252 24622
rect 21196 24518 21252 24556
rect 21420 23380 21476 24782
rect 21644 24612 21700 24622
rect 21644 24162 21700 24556
rect 21980 24388 22036 26126
rect 23100 26180 23156 26190
rect 23100 26178 23268 26180
rect 23100 26126 23102 26178
rect 23154 26126 23268 26178
rect 23100 26124 23268 26126
rect 23100 26114 23156 26124
rect 21980 24322 22036 24332
rect 22092 26068 22148 26078
rect 21644 24110 21646 24162
rect 21698 24110 21700 24162
rect 21644 24098 21700 24110
rect 21868 24276 21924 24286
rect 21868 23938 21924 24220
rect 22092 24050 22148 26012
rect 22672 25900 22936 25910
rect 22728 25844 22776 25900
rect 22832 25844 22880 25900
rect 22672 25834 22936 25844
rect 23100 25844 23156 25854
rect 23100 25506 23156 25788
rect 23100 25454 23102 25506
rect 23154 25454 23156 25506
rect 23100 25442 23156 25454
rect 23212 25284 23268 26124
rect 23436 26178 23492 26190
rect 23436 26126 23438 26178
rect 23490 26126 23492 26178
rect 23100 25228 23268 25284
rect 23324 25282 23380 25294
rect 23324 25230 23326 25282
rect 23378 25230 23380 25282
rect 22652 24834 22708 24846
rect 22652 24782 22654 24834
rect 22706 24782 22708 24834
rect 22540 24724 22596 24734
rect 22092 23998 22094 24050
rect 22146 23998 22148 24050
rect 22092 23986 22148 23998
rect 22204 24612 22260 24622
rect 22204 24498 22260 24556
rect 22204 24446 22206 24498
rect 22258 24446 22260 24498
rect 22204 24164 22260 24446
rect 22316 24610 22372 24622
rect 22316 24558 22318 24610
rect 22370 24558 22372 24610
rect 22316 24276 22372 24558
rect 22316 24210 22372 24220
rect 22428 24388 22484 24398
rect 22204 24052 22260 24108
rect 22204 23996 22372 24052
rect 21868 23886 21870 23938
rect 21922 23886 21924 23938
rect 21868 23492 21924 23886
rect 21868 23426 21924 23436
rect 21980 23828 22036 23838
rect 21420 23314 21476 23324
rect 21532 23268 21588 23278
rect 21588 23212 21700 23268
rect 21532 23202 21588 23212
rect 21084 22990 21086 23042
rect 21138 22990 21140 23042
rect 21084 22978 21140 22990
rect 20860 22642 20916 22652
rect 21532 22370 21588 22382
rect 21532 22318 21534 22370
rect 21586 22318 21588 22370
rect 20748 22258 20804 22270
rect 20748 22206 20750 22258
rect 20802 22206 20804 22258
rect 20748 21812 20804 22206
rect 20748 21746 20804 21756
rect 20860 22148 20916 22158
rect 20860 21586 20916 22092
rect 21532 21812 21588 22318
rect 20860 21534 20862 21586
rect 20914 21534 20916 21586
rect 20860 21522 20916 21534
rect 21420 21700 21476 21710
rect 20636 21476 20692 21486
rect 20636 20802 20692 21420
rect 21420 21362 21476 21644
rect 21420 21310 21422 21362
rect 21474 21310 21476 21362
rect 21420 21298 21476 21310
rect 20636 20750 20638 20802
rect 20690 20750 20692 20802
rect 20636 20738 20692 20750
rect 20748 20804 20804 20814
rect 20748 20710 20804 20748
rect 21532 20802 21588 21756
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21532 20738 21588 20750
rect 20524 20178 20580 20188
rect 21420 20692 21476 20702
rect 21308 20020 21364 20030
rect 21308 19926 21364 19964
rect 19964 17836 20244 17892
rect 20188 17778 20244 17836
rect 20412 17826 20468 17836
rect 20524 19908 20580 19918
rect 20188 17726 20190 17778
rect 20242 17726 20244 17778
rect 20188 17714 20244 17726
rect 19740 16678 19796 16716
rect 20300 17666 20356 17678
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20076 16100 20132 16110
rect 20076 16006 20132 16044
rect 19628 15092 19796 15148
rect 19404 14578 19460 14588
rect 19628 14532 19684 14542
rect 19068 13972 19124 13982
rect 19124 13916 19236 13972
rect 19068 13906 19124 13916
rect 18956 13746 19012 13758
rect 18956 13694 18958 13746
rect 19010 13694 19012 13746
rect 18956 13634 19012 13694
rect 18956 13582 18958 13634
rect 19010 13582 19012 13634
rect 18956 13570 19012 13582
rect 19180 12404 19236 13916
rect 19628 13186 19684 14476
rect 19628 13134 19630 13186
rect 19682 13134 19684 13186
rect 19628 13122 19684 13134
rect 19740 14418 19796 15092
rect 20300 14868 20356 17614
rect 20524 17554 20580 19852
rect 21084 19906 21140 19918
rect 21084 19854 21086 19906
rect 21138 19854 21140 19906
rect 21084 19572 21140 19854
rect 21084 19506 21140 19516
rect 21420 19346 21476 20636
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 21420 19282 21476 19294
rect 21532 20468 21588 20478
rect 21532 19234 21588 20412
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21532 19170 21588 19182
rect 20636 19010 20692 19022
rect 20636 18958 20638 19010
rect 20690 18958 20692 19010
rect 20636 18900 20692 18958
rect 20636 18834 20692 18844
rect 20748 18452 20804 18462
rect 20748 18358 20804 18396
rect 21308 18452 21364 18462
rect 20524 17502 20526 17554
rect 20578 17502 20580 17554
rect 20524 17490 20580 17502
rect 20972 18338 21028 18350
rect 20972 18286 20974 18338
rect 21026 18286 21028 18338
rect 20412 16884 20468 16894
rect 20412 16790 20468 16828
rect 20748 16548 20804 16558
rect 20300 14802 20356 14812
rect 20412 16324 20468 16334
rect 19740 14366 19742 14418
rect 19794 14366 19796 14418
rect 19292 13076 19348 13086
rect 19292 12982 19348 13020
rect 19740 13076 19796 14366
rect 19740 13010 19796 13020
rect 20188 12964 20244 12974
rect 20412 12964 20468 16268
rect 20636 13076 20692 13086
rect 20636 12982 20692 13020
rect 20244 12908 20468 12964
rect 20188 12870 20244 12908
rect 19964 12740 20020 12750
rect 19628 12404 19684 12414
rect 18900 12348 19012 12404
rect 18844 12310 18900 12348
rect 18396 12238 18398 12290
rect 18450 12238 18452 12290
rect 18396 12226 18452 12238
rect 18956 12068 19012 12348
rect 19068 12402 19684 12404
rect 19068 12350 19630 12402
rect 19682 12350 19684 12402
rect 19068 12348 19684 12350
rect 19068 12290 19124 12348
rect 19628 12338 19684 12348
rect 19068 12238 19070 12290
rect 19122 12238 19124 12290
rect 19068 12226 19124 12238
rect 19180 12180 19236 12190
rect 19180 12086 19236 12124
rect 18956 12012 19124 12068
rect 18844 11844 18900 11854
rect 18844 11508 18900 11788
rect 19068 11788 19124 12012
rect 19068 11732 19460 11788
rect 18956 11508 19012 11518
rect 18844 11506 19348 11508
rect 18844 11454 18958 11506
rect 19010 11454 19348 11506
rect 18844 11452 19348 11454
rect 18956 11442 19012 11452
rect 19292 11394 19348 11452
rect 19292 11342 19294 11394
rect 19346 11342 19348 11394
rect 19292 11330 19348 11342
rect 18284 10658 18340 10668
rect 19292 10724 19348 10734
rect 19292 10630 19348 10668
rect 17668 10556 17780 10612
rect 17612 10518 17668 10556
rect 17052 10434 17108 10444
rect 16268 9538 16324 9548
rect 16716 10386 16772 10398
rect 16716 10334 16718 10386
rect 16770 10334 16772 10386
rect 16716 8932 16772 10334
rect 16828 10386 16884 10398
rect 16828 10334 16830 10386
rect 16882 10334 16884 10386
rect 16828 9828 16884 10334
rect 17836 10388 17892 10398
rect 17836 10294 17892 10332
rect 18060 10386 18116 10398
rect 18060 10334 18062 10386
rect 18114 10334 18116 10386
rect 16828 9762 16884 9772
rect 18060 9828 18116 10334
rect 18508 10386 18564 10398
rect 18508 10334 18510 10386
rect 18562 10334 18564 10386
rect 18060 9762 18116 9772
rect 18284 9940 18340 9950
rect 17836 9716 17892 9726
rect 17836 9622 17892 9660
rect 18284 9380 18340 9884
rect 18060 9324 18340 9380
rect 17724 9156 17780 9166
rect 18060 9156 18116 9324
rect 18508 9268 18564 10334
rect 18956 9940 19012 9950
rect 18956 9826 19012 9884
rect 18956 9774 18958 9826
rect 19010 9774 19012 9826
rect 18956 9762 19012 9774
rect 19180 9828 19236 9838
rect 18844 9716 18900 9726
rect 18844 9622 18900 9660
rect 17780 9154 18116 9156
rect 17780 9102 18062 9154
rect 18114 9102 18116 9154
rect 17780 9100 18116 9102
rect 17724 9062 17780 9100
rect 18060 9090 18116 9100
rect 18172 9212 18564 9268
rect 16716 8866 16772 8876
rect 17836 8932 17892 8942
rect 15932 8530 15988 8540
rect 16380 8596 16436 8606
rect 15596 8146 15652 8204
rect 15596 8094 15598 8146
rect 15650 8094 15652 8146
rect 15596 8082 15652 8094
rect 15708 8148 15764 8158
rect 15708 8054 15764 8092
rect 15260 7982 15262 8034
rect 15314 7982 15316 8034
rect 15260 6804 15316 7982
rect 15372 8034 15428 8046
rect 15372 7982 15374 8034
rect 15426 7982 15428 8034
rect 15372 7474 15428 7982
rect 15518 7868 15782 7878
rect 15574 7812 15622 7868
rect 15678 7812 15726 7868
rect 15518 7802 15782 7812
rect 15372 7422 15374 7474
rect 15426 7422 15428 7474
rect 15372 7410 15428 7422
rect 15932 7364 15988 7374
rect 15932 7362 16100 7364
rect 15932 7310 15934 7362
rect 15986 7310 16100 7362
rect 15932 7308 16100 7310
rect 15932 7298 15988 7308
rect 15932 7140 15988 7150
rect 15596 6804 15652 6814
rect 15260 6802 15652 6804
rect 15260 6750 15598 6802
rect 15650 6750 15652 6802
rect 15260 6748 15652 6750
rect 15596 6738 15652 6748
rect 15932 6690 15988 7084
rect 16044 6804 16100 7308
rect 16044 6738 16100 6748
rect 16156 6914 16212 6926
rect 16156 6862 16158 6914
rect 16210 6862 16212 6914
rect 15932 6638 15934 6690
rect 15986 6638 15988 6690
rect 15932 6626 15988 6638
rect 15518 6300 15782 6310
rect 15574 6244 15622 6300
rect 15678 6244 15726 6300
rect 15518 6234 15782 6244
rect 14812 5954 14868 5964
rect 15596 5460 15652 5470
rect 13356 5180 13636 5236
rect 13580 5124 13636 5180
rect 13804 5234 13860 5246
rect 13804 5182 13806 5234
rect 13858 5182 13860 5234
rect 13804 5124 13860 5182
rect 13580 5122 13748 5124
rect 13580 5070 13582 5122
rect 13634 5070 13748 5122
rect 13580 5068 13748 5070
rect 13580 5058 13636 5068
rect 12908 5012 12964 5022
rect 12796 4898 12852 4910
rect 12796 4846 12798 4898
rect 12850 4846 12852 4898
rect 12796 4564 12852 4846
rect 12796 4498 12852 4508
rect 11788 4386 11844 4396
rect 12908 4450 12964 4956
rect 13468 4564 13524 4574
rect 13468 4470 13524 4508
rect 12908 4398 12910 4450
rect 12962 4398 12964 4450
rect 12908 4386 12964 4398
rect 11004 4286 11006 4338
rect 11058 4286 11060 4338
rect 11004 4274 11060 4286
rect 12012 4340 12068 4350
rect 12012 4246 12068 4284
rect 12460 4340 12516 4350
rect 12460 4246 12516 4284
rect 13244 4338 13300 4350
rect 13244 4286 13246 4338
rect 13298 4286 13300 4338
rect 11452 4228 11508 4238
rect 11452 4134 11508 4172
rect 13132 4228 13188 4238
rect 8365 3948 8629 3958
rect 8421 3892 8469 3948
rect 8525 3892 8573 3948
rect 8365 3882 8629 3892
rect 6972 3666 7252 3668
rect 6972 3614 7198 3666
rect 7250 3614 7252 3666
rect 6972 3612 7252 3614
rect 6972 3556 7028 3612
rect 7196 3602 7252 3612
rect 6524 3502 6526 3554
rect 6578 3502 6580 3554
rect 6524 3490 6580 3502
rect 6748 3500 7028 3556
rect 13132 3554 13188 4172
rect 13244 3666 13300 4286
rect 13356 4340 13412 4350
rect 13356 4246 13412 4284
rect 13692 4116 13748 5068
rect 13804 4338 13860 5068
rect 15596 5122 15652 5404
rect 15596 5070 15598 5122
rect 15650 5070 15652 5122
rect 15596 5058 15652 5070
rect 16156 5348 16212 6862
rect 16380 6690 16436 8540
rect 17836 7474 17892 8876
rect 18172 7924 18228 9212
rect 19180 9154 19236 9772
rect 19180 9102 19182 9154
rect 19234 9102 19236 9154
rect 19180 9090 19236 9102
rect 18284 9042 18340 9054
rect 18284 8990 18286 9042
rect 18338 8990 18340 9042
rect 18284 8484 18340 8990
rect 18284 8418 18340 8428
rect 18508 9042 18564 9054
rect 18508 8990 18510 9042
rect 18562 8990 18564 9042
rect 17836 7422 17838 7474
rect 17890 7422 17892 7474
rect 17836 7410 17892 7422
rect 18060 7868 18228 7924
rect 18060 7476 18116 7868
rect 18172 7700 18228 7710
rect 18172 7698 18452 7700
rect 18172 7646 18174 7698
rect 18226 7646 18452 7698
rect 18172 7644 18452 7646
rect 18172 7634 18228 7644
rect 18172 7476 18228 7486
rect 18060 7474 18340 7476
rect 18060 7422 18174 7474
rect 18226 7422 18340 7474
rect 18060 7420 18340 7422
rect 18172 7410 18228 7420
rect 17500 6804 17556 6814
rect 17500 6710 17556 6748
rect 18172 6804 18228 6814
rect 16380 6638 16382 6690
rect 16434 6638 16436 6690
rect 16380 6626 16436 6638
rect 17388 6692 17444 6702
rect 17388 6598 17444 6636
rect 18172 6690 18228 6748
rect 18172 6638 18174 6690
rect 18226 6638 18228 6690
rect 18172 6626 18228 6638
rect 18284 6692 18340 7420
rect 18284 6626 18340 6636
rect 18060 6578 18116 6590
rect 18060 6526 18062 6578
rect 18114 6526 18116 6578
rect 18060 6020 18116 6526
rect 18396 6244 18452 7644
rect 18508 7476 18564 8990
rect 18732 9044 18788 9054
rect 19068 9044 19124 9054
rect 18732 9042 19124 9044
rect 18732 8990 18734 9042
rect 18786 8990 19070 9042
rect 19122 8990 19124 9042
rect 18732 8988 19124 8990
rect 18732 8978 18788 8988
rect 19068 8978 19124 8988
rect 18508 7382 18564 7420
rect 18620 8930 18676 8942
rect 18620 8878 18622 8930
rect 18674 8878 18676 8930
rect 18620 6804 18676 8878
rect 19404 8708 19460 11732
rect 19628 11284 19684 11294
rect 19628 11282 19908 11284
rect 19628 11230 19630 11282
rect 19682 11230 19908 11282
rect 19628 11228 19908 11230
rect 19628 11218 19684 11228
rect 19516 11170 19572 11182
rect 19516 11118 19518 11170
rect 19570 11118 19572 11170
rect 19516 10836 19572 11118
rect 19516 10780 19684 10836
rect 19628 8932 19684 10780
rect 19852 10388 19908 11228
rect 19964 10724 20020 12684
rect 20748 11396 20804 16492
rect 20972 15988 21028 18286
rect 21308 16322 21364 18396
rect 21532 18338 21588 18350
rect 21532 18286 21534 18338
rect 21586 18286 21588 18338
rect 21532 17668 21588 18286
rect 21532 17602 21588 17612
rect 21308 16270 21310 16322
rect 21362 16270 21364 16322
rect 21308 16258 21364 16270
rect 21420 17556 21476 17566
rect 20972 15922 21028 15932
rect 21084 16212 21140 16222
rect 21084 15148 21140 16156
rect 21420 16100 21476 17500
rect 21644 16322 21700 23212
rect 21980 23156 22036 23772
rect 22204 23828 22260 23838
rect 22204 23734 22260 23772
rect 22316 23604 22372 23996
rect 22428 23826 22484 24332
rect 22428 23774 22430 23826
rect 22482 23774 22484 23826
rect 22428 23716 22484 23774
rect 22540 23828 22596 24668
rect 22652 24500 22708 24782
rect 22652 24434 22708 24444
rect 22672 24332 22936 24342
rect 22728 24276 22776 24332
rect 22832 24276 22880 24332
rect 22672 24266 22936 24276
rect 22540 23762 22596 23772
rect 22764 24164 22820 24174
rect 22764 23826 22820 24108
rect 22764 23774 22766 23826
rect 22818 23774 22820 23826
rect 22764 23762 22820 23774
rect 22428 23650 22484 23660
rect 21868 23154 22036 23156
rect 21868 23102 21982 23154
rect 22034 23102 22036 23154
rect 21868 23100 22036 23102
rect 21868 22596 21924 23100
rect 21980 23090 22036 23100
rect 22204 23548 22372 23604
rect 22540 23604 22596 23614
rect 21868 20130 21924 22540
rect 22204 22482 22260 23548
rect 22316 23380 22372 23390
rect 22316 23286 22372 23324
rect 22540 23378 22596 23548
rect 22540 23326 22542 23378
rect 22594 23326 22596 23378
rect 22540 23314 22596 23326
rect 22652 23156 22708 23166
rect 23100 23156 23156 25228
rect 23324 23492 23380 25230
rect 23436 24836 23492 26126
rect 24668 26180 24724 26190
rect 23660 26068 23716 26078
rect 23660 25974 23716 26012
rect 23996 26068 24052 26078
rect 23996 25974 24052 26012
rect 24668 25506 24724 26124
rect 25452 26180 25508 26190
rect 25452 26086 25508 26124
rect 26012 26180 26068 26190
rect 26460 26180 26516 26190
rect 26012 26178 26516 26180
rect 26012 26126 26014 26178
rect 26066 26126 26462 26178
rect 26514 26126 26516 26178
rect 26012 26124 26516 26126
rect 25228 26068 25284 26078
rect 25228 25732 25284 26012
rect 26012 25844 26068 26124
rect 26012 25778 26068 25788
rect 26236 25844 26292 25854
rect 25228 25730 25844 25732
rect 25228 25678 25230 25730
rect 25282 25678 25844 25730
rect 25228 25676 25844 25678
rect 25228 25666 25284 25676
rect 24668 25454 24670 25506
rect 24722 25454 24724 25506
rect 24668 25442 24724 25454
rect 23436 24770 23492 24780
rect 23884 25394 23940 25406
rect 23884 25342 23886 25394
rect 23938 25342 23940 25394
rect 23884 23940 23940 25342
rect 24444 25394 24500 25406
rect 25564 25396 25620 25406
rect 24444 25342 24446 25394
rect 24498 25342 24500 25394
rect 24444 24500 24500 25342
rect 25228 25394 25620 25396
rect 25228 25342 25566 25394
rect 25618 25342 25620 25394
rect 25228 25340 25620 25342
rect 24668 24836 24724 24846
rect 24668 24742 24724 24780
rect 24332 23940 24388 23950
rect 23884 23938 24388 23940
rect 23884 23886 24334 23938
rect 24386 23886 24388 23938
rect 23884 23884 24388 23886
rect 24332 23874 24388 23884
rect 24444 23716 24500 24444
rect 24780 23938 24836 23950
rect 24780 23886 24782 23938
rect 24834 23886 24836 23938
rect 24780 23828 24836 23886
rect 24780 23762 24836 23772
rect 23324 23426 23380 23436
rect 24220 23660 24500 23716
rect 23324 23156 23380 23166
rect 22652 23154 23156 23156
rect 22652 23102 22654 23154
rect 22706 23102 23156 23154
rect 22652 23100 23156 23102
rect 23212 23154 23380 23156
rect 23212 23102 23326 23154
rect 23378 23102 23380 23154
rect 23212 23100 23380 23102
rect 22652 23044 22708 23100
rect 22204 22430 22206 22482
rect 22258 22430 22260 22482
rect 22204 22372 22260 22430
rect 22204 22306 22260 22316
rect 22316 22988 22708 23044
rect 22204 21588 22260 21598
rect 22316 21588 22372 22988
rect 22672 22764 22936 22774
rect 22728 22708 22776 22764
rect 22832 22708 22880 22764
rect 22672 22698 22936 22708
rect 22988 22596 23044 22606
rect 22988 22370 23044 22540
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 22306 23044 22318
rect 22428 22260 22484 22270
rect 22540 22260 22596 22270
rect 22428 22258 22540 22260
rect 22428 22206 22430 22258
rect 22482 22206 22540 22258
rect 22428 22204 22540 22206
rect 22428 22194 22484 22204
rect 22260 21532 22372 21588
rect 22428 22036 22484 22046
rect 22204 21522 22260 21532
rect 22428 20468 22484 21980
rect 22540 21588 22596 22204
rect 22764 22148 22820 22158
rect 22764 22054 22820 22092
rect 23212 21924 23268 23100
rect 23324 23090 23380 23100
rect 23884 23156 23940 23166
rect 23884 23062 23940 23100
rect 22764 21868 23268 21924
rect 23436 23042 23492 23054
rect 23436 22990 23438 23042
rect 23490 22990 23492 23042
rect 22764 21810 22820 21868
rect 22764 21758 22766 21810
rect 22818 21758 22820 21810
rect 22764 21746 22820 21758
rect 23100 21588 23156 21598
rect 22540 21586 23156 21588
rect 22540 21534 23102 21586
rect 23154 21534 23156 21586
rect 22540 21532 23156 21534
rect 23100 21522 23156 21532
rect 22672 21196 22936 21206
rect 22728 21140 22776 21196
rect 22832 21140 22880 21196
rect 22672 21130 22936 21140
rect 22540 20804 22596 20814
rect 22540 20690 22596 20748
rect 23324 20804 23380 20814
rect 23324 20710 23380 20748
rect 22540 20638 22542 20690
rect 22594 20638 22596 20690
rect 22540 20626 22596 20638
rect 22652 20580 22708 20590
rect 22652 20486 22708 20524
rect 22428 20412 22596 20468
rect 22540 20244 22596 20412
rect 22764 20244 22820 20254
rect 22540 20242 22820 20244
rect 22540 20190 22766 20242
rect 22818 20190 22820 20242
rect 22540 20188 22820 20190
rect 22764 20178 22820 20188
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 19908 21924 20078
rect 23324 20132 23380 20142
rect 23436 20132 23492 22990
rect 23548 22372 23604 22382
rect 23548 22260 23604 22316
rect 23548 22258 23716 22260
rect 23548 22206 23550 22258
rect 23602 22206 23716 22258
rect 23548 22204 23716 22206
rect 23548 22194 23604 22204
rect 23660 21698 23716 22204
rect 23660 21646 23662 21698
rect 23714 21646 23716 21698
rect 23660 21634 23716 21646
rect 23996 22258 24052 22270
rect 23996 22206 23998 22258
rect 24050 22206 24052 22258
rect 23884 21588 23940 21598
rect 23884 21494 23940 21532
rect 23996 21252 24052 22206
rect 24220 21476 24276 23660
rect 24444 23492 24500 23502
rect 24444 23266 24500 23436
rect 24556 23380 24612 23390
rect 25228 23380 25284 25340
rect 25564 25330 25620 25340
rect 25564 24946 25620 24958
rect 25564 24894 25566 24946
rect 25618 24894 25620 24946
rect 25340 24500 25396 24510
rect 25340 23826 25396 24444
rect 25340 23774 25342 23826
rect 25394 23774 25396 23826
rect 25340 23762 25396 23774
rect 24556 23286 24612 23324
rect 25004 23324 25284 23380
rect 24444 23214 24446 23266
rect 24498 23214 24500 23266
rect 24444 23202 24500 23214
rect 24780 23154 24836 23166
rect 24780 23102 24782 23154
rect 24834 23102 24836 23154
rect 24668 22596 24724 22606
rect 24668 22502 24724 22540
rect 24332 22370 24388 22382
rect 24332 22318 24334 22370
rect 24386 22318 24388 22370
rect 24332 22260 24388 22318
rect 24332 22194 24388 22204
rect 24556 21698 24612 21710
rect 24556 21646 24558 21698
rect 24610 21646 24612 21698
rect 24332 21476 24388 21486
rect 24220 21474 24388 21476
rect 24220 21422 24334 21474
rect 24386 21422 24388 21474
rect 24220 21420 24388 21422
rect 24332 21410 24388 21420
rect 23996 21186 24052 21196
rect 24556 21252 24612 21646
rect 24556 21186 24612 21196
rect 24668 21362 24724 21374
rect 24668 21310 24670 21362
rect 24722 21310 24724 21362
rect 23324 20130 23492 20132
rect 23324 20078 23326 20130
rect 23378 20078 23492 20130
rect 23324 20076 23492 20078
rect 23660 21026 23716 21038
rect 23660 20974 23662 21026
rect 23714 20974 23716 21026
rect 23324 20066 23380 20076
rect 21868 19842 21924 19852
rect 23660 19794 23716 20974
rect 23996 20802 24052 20814
rect 23996 20750 23998 20802
rect 24050 20750 24052 20802
rect 23996 20132 24052 20750
rect 24220 20132 24276 20142
rect 23996 20130 24276 20132
rect 23996 20078 24222 20130
rect 24274 20078 24276 20130
rect 23996 20076 24276 20078
rect 23660 19742 23662 19794
rect 23714 19742 23716 19794
rect 22672 19628 22936 19638
rect 22728 19572 22776 19628
rect 22832 19572 22880 19628
rect 22672 19562 22936 19572
rect 23548 19572 23604 19582
rect 23100 19292 23380 19348
rect 22204 19012 22260 19022
rect 22092 18564 22148 18574
rect 21868 17892 21924 17902
rect 21756 17556 21812 17566
rect 21868 17556 21924 17836
rect 21756 17554 21924 17556
rect 21756 17502 21758 17554
rect 21810 17502 21924 17554
rect 21756 17500 21924 17502
rect 21756 17490 21812 17500
rect 21644 16270 21646 16322
rect 21698 16270 21700 16322
rect 21644 16258 21700 16270
rect 21532 16100 21588 16110
rect 21420 16044 21532 16100
rect 21532 15986 21588 16044
rect 21532 15934 21534 15986
rect 21586 15934 21588 15986
rect 21532 15922 21588 15934
rect 21980 15988 22036 15998
rect 21980 15894 22036 15932
rect 21532 15314 21588 15326
rect 21532 15262 21534 15314
rect 21586 15262 21588 15314
rect 21084 15092 21364 15148
rect 21196 13860 21252 13870
rect 21084 13748 21140 13758
rect 21084 13634 21140 13692
rect 21196 13746 21252 13804
rect 21196 13694 21198 13746
rect 21250 13694 21252 13746
rect 21196 13682 21252 13694
rect 21084 13582 21086 13634
rect 21138 13582 21140 13634
rect 21084 13570 21140 13582
rect 21308 11396 21364 15092
rect 21532 14644 21588 15262
rect 22092 15202 22148 18508
rect 22204 18226 22260 18956
rect 22764 19010 22820 19022
rect 22764 18958 22766 19010
rect 22818 18958 22820 19010
rect 22540 18564 22596 18574
rect 22540 18450 22596 18508
rect 22540 18398 22542 18450
rect 22594 18398 22596 18450
rect 22540 18386 22596 18398
rect 22204 18174 22206 18226
rect 22258 18174 22260 18226
rect 22204 18162 22260 18174
rect 22316 18338 22372 18350
rect 22316 18286 22318 18338
rect 22370 18286 22372 18338
rect 22316 16996 22372 18286
rect 22764 18340 22820 18958
rect 22764 18274 22820 18284
rect 23100 18562 23156 19292
rect 23324 19234 23380 19292
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 19170 23380 19182
rect 23100 18510 23102 18562
rect 23154 18510 23156 18562
rect 22672 18060 22936 18070
rect 22728 18004 22776 18060
rect 22832 18004 22880 18060
rect 22672 17994 22936 18004
rect 23100 17892 23156 18510
rect 23100 17826 23156 17836
rect 23212 19122 23268 19134
rect 23212 19070 23214 19122
rect 23266 19070 23268 19122
rect 23212 19012 23268 19070
rect 23212 17556 23268 18956
rect 23436 18564 23492 18574
rect 23548 18564 23604 19516
rect 23492 18508 23604 18564
rect 23212 17490 23268 17500
rect 23324 18340 23380 18350
rect 23324 17220 23380 18284
rect 23436 17666 23492 18508
rect 23436 17614 23438 17666
rect 23490 17614 23492 17666
rect 23436 17602 23492 17614
rect 23548 17220 23604 17230
rect 23324 17164 23492 17220
rect 22428 16996 22484 17006
rect 22316 16940 22428 16996
rect 22428 16770 22484 16940
rect 22764 16994 22820 17006
rect 22764 16942 22766 16994
rect 22818 16942 22820 16994
rect 22428 16718 22430 16770
rect 22482 16718 22484 16770
rect 22428 16706 22484 16718
rect 22540 16882 22596 16894
rect 22540 16830 22542 16882
rect 22594 16830 22596 16882
rect 22204 16100 22260 16110
rect 22204 16006 22260 16044
rect 22540 16100 22596 16830
rect 22764 16660 22820 16942
rect 23324 16996 23380 17006
rect 23324 16902 23380 16940
rect 23212 16772 23268 16782
rect 23436 16772 23492 17164
rect 22764 16604 23156 16660
rect 22672 16492 22936 16502
rect 22728 16436 22776 16492
rect 22832 16436 22880 16492
rect 22672 16426 22936 16436
rect 22764 16100 22820 16110
rect 22540 16098 22820 16100
rect 22540 16046 22766 16098
rect 22818 16046 22820 16098
rect 22540 16044 22820 16046
rect 22316 15876 22372 15886
rect 22316 15426 22372 15820
rect 22316 15374 22318 15426
rect 22370 15374 22372 15426
rect 22316 15362 22372 15374
rect 22092 15150 22094 15202
rect 22146 15150 22148 15202
rect 22092 15138 22148 15150
rect 22428 15204 22484 15214
rect 21532 13522 21588 14588
rect 21868 14642 21924 14654
rect 21868 14590 21870 14642
rect 21922 14590 21924 14642
rect 21644 14530 21700 14542
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21644 13860 21700 14478
rect 21868 14532 21924 14590
rect 22428 14642 22484 15148
rect 22428 14590 22430 14642
rect 22482 14590 22484 14642
rect 22428 14578 22484 14590
rect 21868 14466 21924 14476
rect 22540 13970 22596 16044
rect 22764 16034 22820 16044
rect 23100 15538 23156 16604
rect 23212 16100 23268 16716
rect 23212 16006 23268 16044
rect 23324 16716 23492 16772
rect 23548 16882 23604 17164
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 23100 15486 23102 15538
rect 23154 15486 23156 15538
rect 23100 15474 23156 15486
rect 23324 15538 23380 16716
rect 23436 16322 23492 16334
rect 23436 16270 23438 16322
rect 23490 16270 23492 16322
rect 23436 16212 23492 16270
rect 23436 16146 23492 16156
rect 23324 15486 23326 15538
rect 23378 15486 23380 15538
rect 23324 15474 23380 15486
rect 23436 15314 23492 15326
rect 23436 15262 23438 15314
rect 23490 15262 23492 15314
rect 23436 15148 23492 15262
rect 23324 15092 23492 15148
rect 22672 14924 22936 14934
rect 22728 14868 22776 14924
rect 22832 14868 22880 14924
rect 22672 14858 22936 14868
rect 22652 14532 22708 14542
rect 22876 14532 22932 14542
rect 22652 14530 22932 14532
rect 22652 14478 22654 14530
rect 22706 14478 22878 14530
rect 22930 14478 22932 14530
rect 22652 14476 22932 14478
rect 22652 14466 22708 14476
rect 22876 14466 22932 14476
rect 23324 14532 23380 15092
rect 23324 14466 23380 14476
rect 23436 14980 23492 14990
rect 23212 14418 23268 14430
rect 23212 14366 23214 14418
rect 23266 14366 23268 14418
rect 23100 14306 23156 14318
rect 23100 14254 23102 14306
rect 23154 14254 23156 14306
rect 22540 13918 22542 13970
rect 22594 13918 22596 13970
rect 22540 13906 22596 13918
rect 22988 14196 23044 14206
rect 21980 13860 22036 13870
rect 21700 13858 22036 13860
rect 21700 13806 21982 13858
rect 22034 13806 22036 13858
rect 21700 13804 22036 13806
rect 21644 13794 21700 13804
rect 21980 13794 22036 13804
rect 21532 13470 21534 13522
rect 21586 13470 21588 13522
rect 21532 13458 21588 13470
rect 22204 13524 22260 13534
rect 22988 13524 23044 14140
rect 23100 13860 23156 14254
rect 23100 13794 23156 13804
rect 23212 13524 23268 14366
rect 23324 13972 23380 13982
rect 23436 13972 23492 14924
rect 23548 14532 23604 16830
rect 23660 16884 23716 19742
rect 23772 19572 23828 19582
rect 23772 19458 23828 19516
rect 23772 19406 23774 19458
rect 23826 19406 23828 19458
rect 23772 19394 23828 19406
rect 23996 19236 24052 19246
rect 24220 19236 24276 20076
rect 24444 20020 24500 20030
rect 24668 20020 24724 21310
rect 24444 20018 24612 20020
rect 24444 19966 24446 20018
rect 24498 19966 24612 20018
rect 24444 19964 24612 19966
rect 24444 19954 24500 19964
rect 23996 19234 24276 19236
rect 23996 19182 23998 19234
rect 24050 19182 24276 19234
rect 23996 19180 24276 19182
rect 24556 19460 24612 19964
rect 24668 19954 24724 19964
rect 23772 17668 23828 17678
rect 23996 17668 24052 19180
rect 24556 19122 24612 19404
rect 24556 19070 24558 19122
rect 24610 19070 24612 19122
rect 24556 19058 24612 19070
rect 24108 19012 24164 19022
rect 24108 19010 24276 19012
rect 24108 18958 24110 19010
rect 24162 18958 24276 19010
rect 24108 18956 24276 18958
rect 24108 18946 24164 18956
rect 24220 18452 24276 18956
rect 24220 18386 24276 18396
rect 24668 18340 24724 18350
rect 24668 18246 24724 18284
rect 23772 17666 24052 17668
rect 23772 17614 23774 17666
rect 23826 17614 24052 17666
rect 23772 17612 24052 17614
rect 23772 17108 23828 17612
rect 24332 17556 24388 17566
rect 24332 17462 24388 17500
rect 23772 17042 23828 17052
rect 24444 17108 24500 17118
rect 23996 16884 24052 16894
rect 23660 16882 24052 16884
rect 23660 16830 23998 16882
rect 24050 16830 24052 16882
rect 23660 16828 24052 16830
rect 23996 16818 24052 16828
rect 24332 16660 24388 16670
rect 24332 16566 24388 16604
rect 23884 16100 23940 16110
rect 23884 15426 23940 16044
rect 23884 15374 23886 15426
rect 23938 15374 23940 15426
rect 23884 15148 23940 15374
rect 24332 15986 24388 15998
rect 24332 15934 24334 15986
rect 24386 15934 24388 15986
rect 23660 15092 23940 15148
rect 24108 15204 24164 15242
rect 24332 15204 24388 15934
rect 24444 15538 24500 17052
rect 24780 16548 24836 23102
rect 25004 20690 25060 23324
rect 25228 23154 25284 23166
rect 25228 23102 25230 23154
rect 25282 23102 25284 23154
rect 25228 22708 25284 23102
rect 25228 22642 25284 22652
rect 25340 22146 25396 22158
rect 25340 22094 25342 22146
rect 25394 22094 25396 22146
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25004 20638 25006 20690
rect 25058 20638 25060 20690
rect 25004 20626 25060 20638
rect 25116 20802 25172 20814
rect 25116 20750 25118 20802
rect 25170 20750 25172 20802
rect 25116 19346 25172 20750
rect 25228 19572 25284 21534
rect 25340 20804 25396 22094
rect 25340 20738 25396 20748
rect 25228 19506 25284 19516
rect 25340 20580 25396 20590
rect 25116 19294 25118 19346
rect 25170 19294 25172 19346
rect 25116 19282 25172 19294
rect 25004 19234 25060 19246
rect 25004 19182 25006 19234
rect 25058 19182 25060 19234
rect 25004 18676 25060 19182
rect 25004 18610 25060 18620
rect 25228 18452 25284 18462
rect 25228 18358 25284 18396
rect 25340 18004 25396 20524
rect 25564 20018 25620 24894
rect 25676 24722 25732 24734
rect 25676 24670 25678 24722
rect 25730 24670 25732 24722
rect 25676 23380 25732 24670
rect 25788 24610 25844 25676
rect 25788 24558 25790 24610
rect 25842 24558 25844 24610
rect 25788 24546 25844 24558
rect 26124 25508 26180 25518
rect 26236 25508 26292 25788
rect 26460 25620 26516 26124
rect 26460 25554 26516 25564
rect 26124 25506 26292 25508
rect 26124 25454 26126 25506
rect 26178 25454 26292 25506
rect 26124 25452 26292 25454
rect 25676 23314 25732 23324
rect 25788 23604 25844 23614
rect 25676 23044 25732 23054
rect 25676 22950 25732 22988
rect 25676 22260 25732 22270
rect 25788 22260 25844 23548
rect 25676 22258 25844 22260
rect 25676 22206 25678 22258
rect 25730 22206 25844 22258
rect 25676 22204 25844 22206
rect 25676 22036 25732 22204
rect 25676 21970 25732 21980
rect 26124 21700 26180 25452
rect 26684 25396 26740 26350
rect 28924 26404 28980 26414
rect 28924 26310 28980 26348
rect 26348 25394 26740 25396
rect 26348 25342 26686 25394
rect 26738 25342 26740 25394
rect 26348 25340 26740 25342
rect 26236 24052 26292 24062
rect 26236 22258 26292 23996
rect 26348 23492 26404 25340
rect 26684 25330 26740 25340
rect 26908 26290 26964 26302
rect 26908 26238 26910 26290
rect 26962 26238 26964 26290
rect 26684 24724 26740 24734
rect 26908 24724 26964 26238
rect 27356 26292 27412 26302
rect 27132 26178 27188 26190
rect 27132 26126 27134 26178
rect 27186 26126 27188 26178
rect 26684 24722 26964 24724
rect 26684 24670 26686 24722
rect 26738 24670 26964 24722
rect 26684 24668 26964 24670
rect 27020 25956 27076 25966
rect 26460 23716 26516 23726
rect 26684 23716 26740 24668
rect 27020 24500 27076 25900
rect 26460 23714 26684 23716
rect 26460 23662 26462 23714
rect 26514 23662 26684 23714
rect 26460 23660 26684 23662
rect 26460 23650 26516 23660
rect 26684 23622 26740 23660
rect 26908 24444 27076 24500
rect 26348 23426 26404 23436
rect 26460 23044 26516 23054
rect 26460 22950 26516 22988
rect 26796 23042 26852 23054
rect 26796 22990 26798 23042
rect 26850 22990 26852 23042
rect 26796 22708 26852 22990
rect 26796 22642 26852 22652
rect 26236 22206 26238 22258
rect 26290 22206 26292 22258
rect 26236 22194 26292 22206
rect 26572 22370 26628 22382
rect 26572 22318 26574 22370
rect 26626 22318 26628 22370
rect 26572 21812 26628 22318
rect 26796 22260 26852 22270
rect 26796 22166 26852 22204
rect 26572 21718 26628 21756
rect 26460 21700 26516 21710
rect 26124 21634 26180 21644
rect 26348 21698 26516 21700
rect 26348 21646 26462 21698
rect 26514 21646 26516 21698
rect 26348 21644 26516 21646
rect 25676 21476 25732 21486
rect 25676 21382 25732 21420
rect 26348 20244 26404 21644
rect 26460 21634 26516 21644
rect 26908 21588 26964 24444
rect 27132 24052 27188 26126
rect 27356 25844 27412 26236
rect 28700 26292 28756 26302
rect 28756 26236 28868 26292
rect 28700 26198 28756 26236
rect 27692 26180 27748 26190
rect 27692 26178 27860 26180
rect 27692 26126 27694 26178
rect 27746 26126 27860 26178
rect 27692 26124 27860 26126
rect 27692 26114 27748 26124
rect 27356 25778 27412 25788
rect 27692 25508 27748 25518
rect 27244 25506 27748 25508
rect 27244 25454 27694 25506
rect 27746 25454 27748 25506
rect 27244 25452 27748 25454
rect 27244 24834 27300 25452
rect 27692 25442 27748 25452
rect 27804 25284 27860 26124
rect 28476 25396 28532 25406
rect 28476 25302 28532 25340
rect 27244 24782 27246 24834
rect 27298 24782 27300 24834
rect 27244 24770 27300 24782
rect 27692 25228 27860 25284
rect 27132 23996 27412 24052
rect 27356 23938 27412 23996
rect 27356 23886 27358 23938
rect 27410 23886 27412 23938
rect 27356 23874 27412 23886
rect 27132 23492 27188 23502
rect 27020 23380 27076 23390
rect 27020 22596 27076 23324
rect 27132 23154 27188 23436
rect 27132 23102 27134 23154
rect 27186 23102 27188 23154
rect 27132 23090 27188 23102
rect 27132 22596 27188 22606
rect 27020 22594 27188 22596
rect 27020 22542 27134 22594
rect 27186 22542 27188 22594
rect 27020 22540 27188 22542
rect 27132 22530 27188 22540
rect 27692 22484 27748 25228
rect 28364 24724 28420 24734
rect 28364 24630 28420 24668
rect 27804 24610 27860 24622
rect 27804 24558 27806 24610
rect 27858 24558 27860 24610
rect 27804 23940 27860 24558
rect 27804 23846 27860 23884
rect 28476 23938 28532 23950
rect 28476 23886 28478 23938
rect 28530 23886 28532 23938
rect 27356 22428 27748 22484
rect 27916 23826 27972 23838
rect 27916 23774 27918 23826
rect 27970 23774 27972 23826
rect 27132 22372 27188 22382
rect 27356 22372 27412 22428
rect 27132 22370 27412 22372
rect 27132 22318 27134 22370
rect 27186 22318 27412 22370
rect 27132 22316 27412 22318
rect 27020 21588 27076 21598
rect 26908 21532 27020 21588
rect 27020 20914 27076 21532
rect 27020 20862 27022 20914
rect 27074 20862 27076 20914
rect 27020 20850 27076 20862
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25564 19954 25620 19966
rect 25900 20020 25956 20030
rect 25900 19926 25956 19964
rect 26236 19460 26292 19470
rect 25900 19348 25956 19358
rect 25564 19346 25956 19348
rect 25564 19294 25902 19346
rect 25954 19294 25956 19346
rect 25564 19292 25956 19294
rect 25564 19234 25620 19292
rect 25900 19282 25956 19292
rect 26124 19348 26180 19358
rect 25564 19182 25566 19234
rect 25618 19182 25620 19234
rect 25564 19170 25620 19182
rect 26012 19124 26068 19134
rect 25900 19122 26068 19124
rect 25900 19070 26014 19122
rect 26066 19070 26068 19122
rect 25900 19068 26068 19070
rect 25900 19012 25956 19068
rect 26012 19058 26068 19068
rect 25900 18946 25956 18956
rect 25900 18676 25956 18686
rect 25340 17938 25396 17948
rect 25564 18562 25620 18574
rect 25564 18510 25566 18562
rect 25618 18510 25620 18562
rect 25564 18340 25620 18510
rect 25340 17444 25396 17454
rect 25340 17350 25396 17388
rect 25564 16996 25620 18284
rect 25900 18338 25956 18620
rect 26124 18450 26180 19292
rect 26236 19124 26292 19404
rect 26236 19058 26292 19068
rect 26348 18900 26404 20188
rect 26572 20690 26628 20702
rect 26572 20638 26574 20690
rect 26626 20638 26628 20690
rect 26572 20132 26628 20638
rect 26572 20066 26628 20076
rect 27020 19346 27076 19358
rect 27020 19294 27022 19346
rect 27074 19294 27076 19346
rect 27020 19124 27076 19294
rect 27020 19058 27076 19068
rect 26124 18398 26126 18450
rect 26178 18398 26180 18450
rect 26124 18386 26180 18398
rect 26236 18844 26404 18900
rect 26460 19012 26516 19022
rect 25900 18286 25902 18338
rect 25954 18286 25956 18338
rect 25900 18274 25956 18286
rect 26236 18116 26292 18844
rect 26460 18788 26516 18956
rect 26348 18732 26516 18788
rect 26908 18900 26964 18910
rect 26348 18674 26404 18732
rect 26348 18622 26350 18674
rect 26402 18622 26404 18674
rect 26348 18610 26404 18622
rect 26908 18674 26964 18844
rect 26908 18622 26910 18674
rect 26962 18622 26964 18674
rect 26908 18610 26964 18622
rect 26460 18564 26516 18574
rect 26572 18564 26628 18574
rect 26460 18562 26572 18564
rect 26460 18510 26462 18562
rect 26514 18510 26572 18562
rect 26460 18508 26572 18510
rect 26460 18498 26516 18508
rect 25564 16930 25620 16940
rect 25900 18060 26292 18116
rect 24780 16482 24836 16492
rect 24556 16100 24612 16138
rect 24556 16034 24612 16044
rect 25452 16100 25508 16110
rect 24444 15486 24446 15538
rect 24498 15486 24500 15538
rect 24444 15474 24500 15486
rect 24556 15876 24612 15886
rect 24164 15148 24388 15204
rect 24556 15148 24612 15820
rect 25228 15314 25284 15326
rect 25228 15262 25230 15314
rect 25282 15262 25284 15314
rect 25228 15148 25284 15262
rect 25452 15314 25508 16044
rect 25452 15262 25454 15314
rect 25506 15262 25508 15314
rect 25452 15250 25508 15262
rect 24108 15138 24164 15148
rect 24444 15092 24612 15148
rect 25116 15092 25284 15148
rect 25900 15148 25956 18060
rect 26460 17780 26516 17790
rect 26236 17666 26292 17678
rect 26236 17614 26238 17666
rect 26290 17614 26292 17666
rect 26012 17556 26068 17566
rect 26012 16882 26068 17500
rect 26012 16830 26014 16882
rect 26066 16830 26068 16882
rect 26012 15876 26068 16830
rect 26236 17444 26292 17614
rect 26236 16882 26292 17388
rect 26460 17108 26516 17724
rect 26460 16994 26516 17052
rect 26460 16942 26462 16994
rect 26514 16942 26516 16994
rect 26460 16930 26516 16942
rect 26236 16830 26238 16882
rect 26290 16830 26292 16882
rect 26236 16818 26292 16830
rect 26348 16884 26404 16894
rect 26348 16790 26404 16828
rect 26124 16436 26180 16446
rect 26124 16098 26180 16380
rect 26124 16046 26126 16098
rect 26178 16046 26180 16098
rect 26124 16034 26180 16046
rect 26572 16098 26628 18508
rect 26908 16658 26964 16670
rect 26908 16606 26910 16658
rect 26962 16606 26964 16658
rect 26908 16212 26964 16606
rect 27020 16658 27076 16670
rect 27020 16606 27022 16658
rect 27074 16606 27076 16658
rect 27020 16436 27076 16606
rect 27132 16548 27188 22316
rect 27692 21588 27748 21598
rect 27468 20018 27524 20030
rect 27468 19966 27470 20018
rect 27522 19966 27524 20018
rect 27468 19348 27524 19966
rect 27468 19282 27524 19292
rect 27692 19234 27748 21532
rect 27692 19182 27694 19234
rect 27746 19182 27748 19234
rect 27692 18900 27748 19182
rect 27692 18834 27748 18844
rect 27356 18452 27412 18462
rect 27356 17332 27412 18396
rect 27916 18340 27972 23774
rect 28028 23266 28084 23278
rect 28028 23214 28030 23266
rect 28082 23214 28084 23266
rect 28028 22708 28084 23214
rect 28028 22642 28084 22652
rect 28252 22260 28308 22270
rect 28252 22258 28420 22260
rect 28252 22206 28254 22258
rect 28306 22206 28420 22258
rect 28252 22204 28420 22206
rect 28252 22194 28308 22204
rect 28252 20802 28308 20814
rect 28252 20750 28254 20802
rect 28306 20750 28308 20802
rect 28252 20692 28308 20750
rect 28252 20626 28308 20636
rect 28364 20690 28420 22204
rect 28476 21476 28532 23886
rect 28588 23940 28644 23950
rect 28588 23044 28644 23884
rect 28700 23716 28756 23726
rect 28700 23266 28756 23660
rect 28700 23214 28702 23266
rect 28754 23214 28756 23266
rect 28700 23202 28756 23214
rect 28588 22988 28756 23044
rect 28588 22708 28644 22718
rect 28588 21698 28644 22652
rect 28588 21646 28590 21698
rect 28642 21646 28644 21698
rect 28588 21634 28644 21646
rect 28700 21586 28756 22988
rect 28812 22932 28868 26236
rect 29484 26290 29540 26302
rect 29484 26238 29486 26290
rect 29538 26238 29540 26290
rect 29372 25620 29428 25630
rect 29148 25564 29372 25620
rect 29148 24834 29204 25564
rect 29372 25526 29428 25564
rect 29148 24782 29150 24834
rect 29202 24782 29204 24834
rect 29148 24770 29204 24782
rect 29484 24724 29540 26238
rect 29596 24948 29652 26852
rect 48748 26850 48804 26862
rect 48748 26798 48750 26850
rect 48802 26798 48804 26850
rect 29825 26684 30089 26694
rect 29881 26628 29929 26684
rect 29985 26628 30033 26684
rect 29825 26618 30089 26628
rect 44132 26684 44396 26694
rect 44188 26628 44236 26684
rect 44292 26628 44340 26684
rect 44132 26618 44396 26628
rect 48748 26514 48804 26798
rect 48748 26462 48750 26514
rect 48802 26462 48804 26514
rect 48748 26450 48804 26462
rect 49084 26850 49140 26862
rect 49084 26798 49086 26850
rect 49138 26798 49140 26850
rect 29932 26404 29988 26414
rect 29932 26178 29988 26348
rect 36092 26404 36148 26414
rect 29932 26126 29934 26178
rect 29986 26126 29988 26178
rect 29820 26066 29876 26078
rect 29820 26014 29822 26066
rect 29874 26014 29876 26066
rect 29820 25620 29876 26014
rect 29932 25620 29988 26126
rect 31276 26292 31332 26302
rect 31164 26066 31220 26078
rect 31164 26014 31166 26066
rect 31218 26014 31220 26066
rect 30044 25620 30100 25630
rect 29932 25618 30100 25620
rect 29932 25566 30046 25618
rect 30098 25566 30100 25618
rect 29932 25564 30100 25566
rect 29820 25554 29876 25564
rect 30044 25284 30100 25564
rect 30156 25508 30212 25518
rect 30156 25506 30996 25508
rect 30156 25454 30158 25506
rect 30210 25454 30996 25506
rect 30156 25452 30996 25454
rect 30156 25442 30212 25452
rect 30044 25228 30212 25284
rect 29825 25116 30089 25126
rect 29881 25060 29929 25116
rect 29985 25060 30033 25116
rect 29825 25050 30089 25060
rect 29596 24882 29652 24892
rect 29596 24724 29652 24734
rect 29484 24668 29596 24724
rect 29148 23938 29204 23950
rect 29148 23886 29150 23938
rect 29202 23886 29204 23938
rect 29148 23604 29204 23886
rect 29260 23828 29316 23838
rect 29260 23734 29316 23772
rect 29148 23538 29204 23548
rect 28924 22932 28980 22942
rect 28812 22876 28924 22932
rect 28924 22866 28980 22876
rect 29596 22370 29652 24668
rect 30156 24722 30212 25228
rect 30604 24948 30660 24958
rect 30156 24670 30158 24722
rect 30210 24670 30212 24722
rect 29596 22318 29598 22370
rect 29650 22318 29652 22370
rect 29596 22306 29652 22318
rect 29708 23714 29764 23726
rect 29708 23662 29710 23714
rect 29762 23662 29764 23714
rect 29708 23156 29764 23662
rect 29825 23548 30089 23558
rect 29881 23492 29929 23548
rect 29985 23492 30033 23548
rect 29825 23482 30089 23492
rect 28700 21534 28702 21586
rect 28754 21534 28756 21586
rect 28700 21522 28756 21534
rect 29708 21586 29764 23100
rect 30156 22370 30212 24670
rect 30492 24724 30548 24734
rect 30492 24630 30548 24668
rect 30604 24050 30660 24892
rect 30940 24610 30996 25452
rect 31164 25172 31220 26014
rect 31164 25106 31220 25116
rect 30940 24558 30942 24610
rect 30994 24558 30996 24610
rect 30940 24546 30996 24558
rect 31052 24836 31108 24846
rect 30604 23998 30606 24050
rect 30658 23998 30660 24050
rect 30604 23986 30660 23998
rect 31052 23938 31108 24780
rect 31276 24724 31332 26236
rect 33068 26290 33124 26302
rect 33068 26238 33070 26290
rect 33122 26238 33124 26290
rect 32284 26178 32340 26190
rect 32284 26126 32286 26178
rect 32338 26126 32340 26178
rect 31948 25956 32004 25966
rect 32284 25956 32340 26126
rect 32004 25900 32340 25956
rect 31948 25890 32004 25900
rect 31612 25620 31668 25630
rect 31388 24948 31444 24958
rect 31388 24854 31444 24892
rect 31388 24724 31444 24734
rect 31276 24668 31388 24724
rect 31388 24658 31444 24668
rect 31052 23886 31054 23938
rect 31106 23886 31108 23938
rect 30380 23492 30436 23502
rect 30380 23154 30436 23436
rect 31052 23380 31108 23886
rect 30380 23102 30382 23154
rect 30434 23102 30436 23154
rect 30380 22932 30436 23102
rect 30828 23154 30884 23166
rect 30828 23102 30830 23154
rect 30882 23102 30884 23154
rect 30492 23044 30548 23054
rect 30492 22950 30548 22988
rect 30380 22820 30436 22876
rect 30380 22764 30548 22820
rect 30156 22318 30158 22370
rect 30210 22318 30212 22370
rect 30156 22306 30212 22318
rect 29825 21980 30089 21990
rect 29881 21924 29929 21980
rect 29985 21924 30033 21980
rect 29825 21914 30089 21924
rect 29708 21534 29710 21586
rect 29762 21534 29764 21586
rect 29708 21522 29764 21534
rect 30380 21812 30436 21822
rect 28476 21410 28532 21420
rect 30156 21474 30212 21486
rect 30156 21422 30158 21474
rect 30210 21422 30212 21474
rect 28364 20638 28366 20690
rect 28418 20638 28420 20690
rect 27916 18274 27972 18284
rect 28028 19124 28084 19134
rect 28364 19124 28420 20638
rect 29148 20802 29204 20814
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 29148 20244 29204 20750
rect 28588 20018 28644 20030
rect 28588 19966 28590 20018
rect 28642 19966 28644 20018
rect 28028 19122 28420 19124
rect 28028 19070 28030 19122
rect 28082 19070 28420 19122
rect 28028 19068 28420 19070
rect 28476 19236 28532 19246
rect 28028 18562 28084 19068
rect 28028 18510 28030 18562
rect 28082 18510 28084 18562
rect 28028 17892 28084 18510
rect 28028 17826 28084 17836
rect 28476 17890 28532 19180
rect 28588 18676 28644 19966
rect 29148 19234 29204 20188
rect 29148 19182 29150 19234
rect 29202 19182 29204 19234
rect 29148 19170 29204 19182
rect 29372 20692 29428 20702
rect 29372 19234 29428 20636
rect 29820 20692 29876 20702
rect 29820 20598 29876 20636
rect 29825 20412 30089 20422
rect 29881 20356 29929 20412
rect 29985 20356 30033 20412
rect 29825 20346 30089 20356
rect 30156 20244 30212 21422
rect 30156 20178 30212 20188
rect 30268 21252 30324 21262
rect 30044 20018 30100 20030
rect 30044 19966 30046 20018
rect 30098 19966 30100 20018
rect 29484 19796 29540 19806
rect 29484 19702 29540 19740
rect 30044 19348 30100 19966
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 28588 18610 28644 18620
rect 28700 18674 28756 18686
rect 28700 18622 28702 18674
rect 28754 18622 28756 18674
rect 28700 18564 28756 18622
rect 28700 18498 28756 18508
rect 28476 17838 28478 17890
rect 28530 17838 28532 17890
rect 28476 17826 28532 17838
rect 29148 18452 29204 18462
rect 29372 18452 29428 19182
rect 29708 19292 30044 19348
rect 29708 18564 29764 19292
rect 30044 19282 30100 19292
rect 30268 19346 30324 21196
rect 30380 20802 30436 21756
rect 30380 20750 30382 20802
rect 30434 20750 30436 20802
rect 30380 20738 30436 20750
rect 30492 20690 30548 22764
rect 30828 22258 30884 23102
rect 31052 23154 31108 23324
rect 31052 23102 31054 23154
rect 31106 23102 31108 23154
rect 31052 23090 31108 23102
rect 31388 23044 31444 23054
rect 30828 22206 30830 22258
rect 30882 22206 30884 22258
rect 30492 20638 30494 20690
rect 30546 20638 30548 20690
rect 30492 20626 30548 20638
rect 30604 20692 30660 20702
rect 30492 20132 30548 20142
rect 30268 19294 30270 19346
rect 30322 19294 30324 19346
rect 30268 19282 30324 19294
rect 30380 20130 30548 20132
rect 30380 20078 30494 20130
rect 30546 20078 30548 20130
rect 30380 20076 30548 20078
rect 29825 18844 30089 18854
rect 29881 18788 29929 18844
rect 29985 18788 30033 18844
rect 29825 18778 30089 18788
rect 29596 18452 29652 18462
rect 29204 18450 29652 18452
rect 29204 18398 29598 18450
rect 29650 18398 29652 18450
rect 29204 18396 29652 18398
rect 28364 17668 28420 17678
rect 28364 17574 28420 17612
rect 27692 17556 27748 17566
rect 27692 17462 27748 17500
rect 27356 17266 27412 17276
rect 28364 17220 28420 17230
rect 27916 17108 27972 17118
rect 27580 17106 27972 17108
rect 27580 17054 27918 17106
rect 27970 17054 27972 17106
rect 27580 17052 27972 17054
rect 27244 16996 27300 17006
rect 27244 16770 27300 16940
rect 27356 16884 27412 16894
rect 27580 16884 27636 17052
rect 27916 17042 27972 17052
rect 27356 16882 27636 16884
rect 27356 16830 27358 16882
rect 27410 16830 27636 16882
rect 27356 16828 27636 16830
rect 27692 16884 27748 16894
rect 27356 16818 27412 16828
rect 27692 16790 27748 16828
rect 28364 16884 28420 17164
rect 28364 16882 28644 16884
rect 28364 16830 28366 16882
rect 28418 16830 28644 16882
rect 28364 16828 28644 16830
rect 28364 16818 28420 16828
rect 27244 16718 27246 16770
rect 27298 16718 27300 16770
rect 27244 16706 27300 16718
rect 27804 16770 27860 16782
rect 27804 16718 27806 16770
rect 27858 16718 27860 16770
rect 27132 16492 27412 16548
rect 27020 16370 27076 16380
rect 27356 16212 27412 16492
rect 26908 16156 27076 16212
rect 26572 16046 26574 16098
rect 26626 16046 26628 16098
rect 26572 16034 26628 16046
rect 26012 15810 26068 15820
rect 26684 15876 26740 15886
rect 26684 15782 26740 15820
rect 26908 15874 26964 15886
rect 26908 15822 26910 15874
rect 26962 15822 26964 15874
rect 26908 15764 26964 15822
rect 26908 15698 26964 15708
rect 27020 15540 27076 16156
rect 27244 16156 27412 16212
rect 27132 16100 27188 16110
rect 27132 16006 27188 16044
rect 27020 15426 27076 15484
rect 27020 15374 27022 15426
rect 27074 15374 27076 15426
rect 27020 15362 27076 15374
rect 27244 15148 27300 16156
rect 27804 16100 27860 16718
rect 27356 16044 27860 16100
rect 27356 15986 27412 16044
rect 27356 15934 27358 15986
rect 27410 15934 27412 15986
rect 27356 15922 27412 15934
rect 27804 15876 27860 16044
rect 27916 16548 27972 16558
rect 27916 16098 27972 16492
rect 28252 16548 28308 16558
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27916 16034 27972 16046
rect 28140 16100 28196 16110
rect 27804 15820 27972 15876
rect 27692 15764 27748 15774
rect 27692 15426 27748 15708
rect 27916 15538 27972 15820
rect 27916 15486 27918 15538
rect 27970 15486 27972 15538
rect 27916 15474 27972 15486
rect 28140 15538 28196 16044
rect 28140 15486 28142 15538
rect 28194 15486 28196 15538
rect 28140 15474 28196 15486
rect 28252 15538 28308 16492
rect 28364 16098 28420 16110
rect 28364 16046 28366 16098
rect 28418 16046 28420 16098
rect 28364 15764 28420 16046
rect 28588 15988 28644 16828
rect 28476 15876 28532 15886
rect 28476 15782 28532 15820
rect 28364 15698 28420 15708
rect 28252 15486 28254 15538
rect 28306 15486 28308 15538
rect 28252 15474 28308 15486
rect 27692 15374 27694 15426
rect 27746 15374 27748 15426
rect 27692 15362 27748 15374
rect 25900 15092 26068 15148
rect 23660 14642 23716 15092
rect 24444 14868 24500 15092
rect 24220 14812 24500 14868
rect 24780 14980 24836 14990
rect 24220 14754 24276 14812
rect 24220 14702 24222 14754
rect 24274 14702 24276 14754
rect 24220 14690 24276 14702
rect 23660 14590 23662 14642
rect 23714 14590 23716 14642
rect 23660 14578 23716 14590
rect 23884 14644 23940 14654
rect 23884 14550 23940 14588
rect 23548 14466 23604 14476
rect 24444 14532 24500 14542
rect 24444 14438 24500 14476
rect 24780 14530 24836 14924
rect 25116 14644 25172 15092
rect 25116 14578 25172 14588
rect 24780 14478 24782 14530
rect 24834 14478 24836 14530
rect 23324 13970 23492 13972
rect 23324 13918 23326 13970
rect 23378 13918 23492 13970
rect 23324 13916 23492 13918
rect 23772 14196 23828 14206
rect 23772 13970 23828 14140
rect 23772 13918 23774 13970
rect 23826 13918 23828 13970
rect 23324 13906 23380 13916
rect 23772 13906 23828 13918
rect 24780 13972 24836 14478
rect 26012 14418 26068 15092
rect 27132 15092 27300 15148
rect 28252 15316 28308 15326
rect 28252 15202 28308 15260
rect 28252 15150 28254 15202
rect 28306 15150 28308 15202
rect 28252 15138 28308 15150
rect 26796 14756 26852 14766
rect 26012 14366 26014 14418
rect 26066 14366 26068 14418
rect 22988 13468 23156 13524
rect 22204 13430 22260 13468
rect 21420 13412 21476 13422
rect 21420 13076 21476 13356
rect 22672 13356 22936 13366
rect 22728 13300 22776 13356
rect 22832 13300 22880 13356
rect 22672 13290 22936 13300
rect 22092 13188 22148 13198
rect 21420 13074 21588 13076
rect 21420 13022 21422 13074
rect 21474 13022 21588 13074
rect 21420 13020 21588 13022
rect 21420 13010 21476 13020
rect 21532 12516 21588 13020
rect 21868 12964 21924 12974
rect 21924 12908 22036 12964
rect 21868 12870 21924 12908
rect 21532 12460 21924 12516
rect 21644 12068 21700 12078
rect 21644 11974 21700 12012
rect 21868 11618 21924 12460
rect 21980 12068 22036 12908
rect 22092 12402 22148 13132
rect 22988 13188 23044 13198
rect 22540 13076 22596 13086
rect 22092 12350 22094 12402
rect 22146 12350 22148 12402
rect 22092 12338 22148 12350
rect 22316 12850 22372 12862
rect 22316 12798 22318 12850
rect 22370 12798 22372 12850
rect 21980 12002 22036 12012
rect 22204 11956 22260 11966
rect 21868 11566 21870 11618
rect 21922 11566 21924 11618
rect 21868 11554 21924 11566
rect 22092 11620 22148 11630
rect 22204 11620 22260 11900
rect 22092 11618 22260 11620
rect 22092 11566 22094 11618
rect 22146 11566 22260 11618
rect 22092 11564 22260 11566
rect 22316 11620 22372 12798
rect 22540 12402 22596 13020
rect 22988 13074 23044 13132
rect 22988 13022 22990 13074
rect 23042 13022 23044 13074
rect 22988 13010 23044 13022
rect 22540 12350 22542 12402
rect 22594 12350 22596 12402
rect 22540 12338 22596 12350
rect 22988 12404 23044 12414
rect 23100 12404 23156 13468
rect 23212 13458 23268 13468
rect 24332 13634 24388 13646
rect 24332 13582 24334 13634
rect 24386 13582 24388 13634
rect 24332 13524 24388 13582
rect 24668 13636 24724 13646
rect 24668 13542 24724 13580
rect 24332 13458 24388 13468
rect 23772 13188 23828 13198
rect 23324 13076 23380 13086
rect 23324 12962 23380 13020
rect 23324 12910 23326 12962
rect 23378 12910 23380 12962
rect 23324 12898 23380 12910
rect 22988 12402 23100 12404
rect 22988 12350 22990 12402
rect 23042 12350 23100 12402
rect 22988 12348 23100 12350
rect 22988 12338 23044 12348
rect 23100 12310 23156 12348
rect 23100 12180 23156 12190
rect 22672 11788 22936 11798
rect 22728 11732 22776 11788
rect 22832 11732 22880 11788
rect 22672 11722 22936 11732
rect 22316 11564 22708 11620
rect 22092 11554 22148 11564
rect 22316 11396 22372 11406
rect 21308 11340 21588 11396
rect 20748 11302 20804 11340
rect 19964 10658 20020 10668
rect 21420 11170 21476 11182
rect 21420 11118 21422 11170
rect 21474 11118 21476 11170
rect 20748 10610 20804 10622
rect 20748 10558 20750 10610
rect 20802 10558 20804 10610
rect 19964 10388 20020 10398
rect 19852 10332 19964 10388
rect 19964 10050 20020 10332
rect 20748 10388 20804 10558
rect 20748 10322 20804 10332
rect 21084 10610 21140 10622
rect 21084 10558 21086 10610
rect 21138 10558 21140 10610
rect 19964 9998 19966 10050
rect 20018 9998 20020 10050
rect 19964 9986 20020 9998
rect 21084 9156 21140 10558
rect 21084 9090 21140 9100
rect 19628 8866 19684 8876
rect 20412 8932 20468 8942
rect 19404 8652 19908 8708
rect 19852 8258 19908 8652
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8194 19908 8206
rect 20188 8370 20244 8382
rect 20188 8318 20190 8370
rect 20242 8318 20244 8370
rect 20188 8260 20244 8318
rect 18620 6738 18676 6748
rect 19068 7476 19124 7486
rect 18508 6692 18564 6702
rect 18508 6598 18564 6636
rect 18396 6188 18564 6244
rect 18396 6020 18452 6030
rect 18060 6018 18452 6020
rect 18060 5966 18398 6018
rect 18450 5966 18452 6018
rect 18060 5964 18452 5966
rect 18396 5954 18452 5964
rect 18508 5908 18564 6188
rect 19068 6132 19124 7420
rect 20188 7476 20244 8204
rect 20188 7382 20244 7420
rect 20412 7474 20468 8876
rect 21308 8932 21364 8942
rect 21308 8370 21364 8876
rect 21308 8318 21310 8370
rect 21362 8318 21364 8370
rect 21308 8306 21364 8318
rect 20524 8148 20580 8158
rect 20524 8054 20580 8092
rect 20412 7422 20414 7474
rect 20466 7422 20468 7474
rect 20412 7410 20468 7422
rect 21084 7476 21140 7486
rect 21084 7382 21140 7420
rect 21420 7028 21476 11118
rect 21532 9268 21588 11340
rect 22316 11302 22372 11340
rect 22540 11282 22596 11294
rect 22540 11230 22542 11282
rect 22594 11230 22596 11282
rect 21644 10724 21700 10734
rect 21644 10630 21700 10668
rect 21868 10722 21924 10734
rect 21868 10670 21870 10722
rect 21922 10670 21924 10722
rect 21868 10388 21924 10670
rect 22428 10724 22484 10734
rect 22428 10610 22484 10668
rect 22428 10558 22430 10610
rect 22482 10558 22484 10610
rect 21868 10322 21924 10332
rect 21980 10386 22036 10398
rect 21980 10334 21982 10386
rect 22034 10334 22036 10386
rect 21980 9380 22036 10334
rect 22428 9828 22484 10558
rect 22540 10612 22596 11230
rect 22652 11284 22708 11564
rect 22988 11284 23044 11294
rect 22652 11282 23044 11284
rect 22652 11230 22990 11282
rect 23042 11230 23044 11282
rect 22652 11228 23044 11230
rect 22988 11060 23044 11228
rect 23100 11284 23156 12124
rect 23324 12178 23380 12190
rect 23548 12180 23604 12190
rect 23324 12126 23326 12178
rect 23378 12126 23380 12178
rect 23324 11394 23380 12126
rect 23324 11342 23326 11394
rect 23378 11342 23380 11394
rect 23324 11330 23380 11342
rect 23436 12178 23604 12180
rect 23436 12126 23550 12178
rect 23602 12126 23604 12178
rect 23436 12124 23604 12126
rect 23436 11956 23492 12124
rect 23548 12114 23604 12124
rect 23100 11218 23156 11228
rect 22988 11004 23268 11060
rect 22876 10612 22932 10622
rect 22540 10610 22932 10612
rect 22540 10558 22878 10610
rect 22930 10558 22932 10610
rect 22540 10556 22932 10558
rect 22876 10388 22932 10556
rect 22876 10322 22932 10332
rect 22672 10220 22936 10230
rect 22728 10164 22776 10220
rect 22832 10164 22880 10220
rect 22672 10154 22936 10164
rect 22652 9828 22708 9838
rect 22428 9826 22708 9828
rect 22428 9774 22654 9826
rect 22706 9774 22708 9826
rect 22428 9772 22708 9774
rect 22652 9762 22708 9772
rect 23212 9714 23268 11004
rect 23212 9662 23214 9714
rect 23266 9662 23268 9714
rect 23212 9650 23268 9662
rect 23324 10610 23380 10622
rect 23324 10558 23326 10610
rect 23378 10558 23380 10610
rect 23324 9828 23380 10558
rect 23436 10386 23492 11900
rect 23772 11394 23828 13132
rect 24780 13074 24836 13916
rect 25900 13972 25956 13982
rect 25900 13878 25956 13916
rect 25340 13748 25396 13758
rect 25340 13654 25396 13692
rect 25228 13634 25284 13646
rect 25228 13582 25230 13634
rect 25282 13582 25284 13634
rect 25228 13188 25284 13582
rect 25228 13122 25284 13132
rect 24780 13022 24782 13074
rect 24834 13022 24836 13074
rect 24780 13010 24836 13022
rect 23772 11342 23774 11394
rect 23826 11342 23828 11394
rect 23772 11060 23828 11342
rect 23996 12404 24052 12414
rect 23996 11396 24052 12348
rect 24668 12404 24724 12414
rect 24668 12310 24724 12348
rect 25564 12404 25620 12414
rect 25564 12178 25620 12348
rect 25564 12126 25566 12178
rect 25618 12126 25620 12178
rect 25564 12114 25620 12126
rect 24108 12068 24164 12078
rect 24108 12066 24276 12068
rect 24108 12014 24110 12066
rect 24162 12014 24276 12066
rect 24108 12012 24276 12014
rect 24108 12002 24164 12012
rect 23996 11394 24164 11396
rect 23996 11342 23998 11394
rect 24050 11342 24164 11394
rect 23996 11340 24164 11342
rect 23996 11330 24052 11340
rect 23772 10994 23828 11004
rect 24108 10834 24164 11340
rect 24108 10782 24110 10834
rect 24162 10782 24164 10834
rect 24108 10770 24164 10782
rect 23436 10334 23438 10386
rect 23490 10334 23492 10386
rect 23436 10322 23492 10334
rect 21980 9324 22260 9380
rect 21644 9268 21700 9278
rect 21532 9266 22036 9268
rect 21532 9214 21646 9266
rect 21698 9214 22036 9266
rect 21532 9212 22036 9214
rect 21644 9202 21700 9212
rect 21980 9044 22036 9212
rect 21980 8950 22036 8988
rect 21532 8260 21588 8270
rect 21532 8166 21588 8204
rect 21868 8260 21924 8270
rect 22204 8260 22260 9324
rect 22540 9156 22596 9166
rect 22540 9062 22596 9100
rect 22672 8652 22936 8662
rect 22728 8596 22776 8652
rect 22832 8596 22880 8652
rect 22672 8586 22936 8596
rect 23324 8484 23380 9772
rect 24108 9602 24164 9614
rect 24108 9550 24110 9602
rect 24162 9550 24164 9602
rect 23660 9042 23716 9054
rect 23660 8990 23662 9042
rect 23714 8990 23716 9042
rect 23660 8484 23716 8990
rect 22876 8428 23380 8484
rect 23436 8428 23716 8484
rect 22316 8260 22372 8270
rect 22204 8258 22372 8260
rect 22204 8206 22318 8258
rect 22370 8206 22372 8258
rect 22204 8204 22372 8206
rect 21868 8166 21924 8204
rect 22316 8194 22372 8204
rect 22876 8258 22932 8428
rect 22876 8206 22878 8258
rect 22930 8206 22932 8258
rect 22876 8194 22932 8206
rect 23436 8260 23492 8428
rect 23436 7924 23492 8204
rect 23436 7858 23492 7868
rect 23884 8146 23940 8158
rect 23884 8094 23886 8146
rect 23938 8094 23940 8146
rect 21308 6972 21476 7028
rect 22672 7084 22936 7094
rect 22728 7028 22776 7084
rect 22832 7028 22880 7084
rect 22672 7018 22936 7028
rect 20524 6804 20580 6814
rect 19068 6018 19124 6076
rect 19292 6132 19348 6142
rect 19292 6130 19572 6132
rect 19292 6078 19294 6130
rect 19346 6078 19572 6130
rect 19292 6076 19572 6078
rect 19292 6066 19348 6076
rect 19068 5966 19070 6018
rect 19122 5966 19124 6018
rect 19068 5954 19124 5966
rect 19516 6020 19572 6076
rect 19516 5964 19684 6020
rect 18508 5842 18564 5852
rect 18844 5908 18900 5918
rect 18844 5814 18900 5852
rect 19404 5906 19460 5918
rect 19404 5854 19406 5906
rect 19458 5854 19460 5906
rect 18508 5684 18564 5694
rect 19404 5684 19460 5854
rect 18508 5682 18676 5684
rect 18508 5630 18510 5682
rect 18562 5630 18676 5682
rect 18508 5628 18676 5630
rect 18508 5618 18564 5628
rect 13804 4286 13806 4338
rect 13858 4286 13860 4338
rect 13804 4274 13860 4286
rect 13916 5010 13972 5022
rect 13916 4958 13918 5010
rect 13970 4958 13972 5010
rect 13916 4340 13972 4958
rect 15820 5012 15876 5022
rect 15820 4918 15876 4956
rect 15518 4732 15782 4742
rect 15574 4676 15622 4732
rect 15678 4676 15726 4732
rect 15518 4666 15782 4676
rect 13916 4274 13972 4284
rect 14476 4450 14532 4462
rect 14476 4398 14478 4450
rect 14530 4398 14532 4450
rect 14476 4340 14532 4398
rect 16156 4450 16212 5292
rect 17948 5460 18004 5470
rect 16380 5124 16436 5134
rect 16380 5030 16436 5068
rect 16716 4898 16772 4910
rect 16716 4846 16718 4898
rect 16770 4846 16772 4898
rect 16716 4676 16772 4846
rect 16716 4610 16772 4620
rect 16156 4398 16158 4450
rect 16210 4398 16212 4450
rect 16156 4386 16212 4398
rect 16380 4452 16436 4462
rect 16380 4358 16436 4396
rect 14476 4274 14532 4284
rect 17948 4338 18004 5404
rect 18620 5348 18676 5628
rect 19068 5628 19460 5684
rect 18956 5348 19012 5358
rect 19068 5348 19124 5628
rect 18620 5346 19124 5348
rect 18620 5294 18958 5346
rect 19010 5294 19124 5346
rect 18620 5292 19124 5294
rect 19180 5460 19236 5470
rect 18956 5282 19012 5292
rect 18732 5012 18788 5022
rect 18060 4452 18116 4462
rect 18060 4358 18116 4396
rect 17948 4286 17950 4338
rect 18002 4286 18004 4338
rect 17948 4274 18004 4286
rect 18732 4338 18788 4956
rect 19180 5010 19236 5404
rect 19292 5236 19348 5246
rect 19292 5234 19572 5236
rect 19292 5182 19294 5234
rect 19346 5182 19572 5234
rect 19292 5180 19572 5182
rect 19292 5170 19348 5180
rect 19180 4958 19182 5010
rect 19234 4958 19236 5010
rect 19180 4946 19236 4958
rect 19516 4450 19572 5180
rect 19628 5012 19684 5964
rect 19628 4946 19684 4956
rect 19740 5460 19796 5470
rect 19516 4398 19518 4450
rect 19570 4398 19572 4450
rect 19516 4386 19572 4398
rect 19740 4450 19796 5404
rect 20188 5122 20244 5134
rect 20188 5070 20190 5122
rect 20242 5070 20244 5122
rect 20188 4676 20244 5070
rect 20524 5122 20580 6748
rect 21308 5908 21364 6972
rect 23884 6916 23940 8094
rect 23884 6850 23940 6860
rect 21420 6804 21476 6814
rect 21420 6018 21476 6748
rect 24108 6692 24164 9550
rect 23660 6690 24164 6692
rect 23660 6638 24110 6690
rect 24162 6638 24164 6690
rect 23660 6636 24164 6638
rect 23324 6468 23380 6478
rect 21756 6132 21812 6142
rect 21420 5966 21422 6018
rect 21474 5966 21476 6018
rect 21420 5954 21476 5966
rect 21532 6130 21812 6132
rect 21532 6078 21758 6130
rect 21810 6078 21812 6130
rect 21532 6076 21812 6078
rect 21308 5842 21364 5852
rect 20524 5070 20526 5122
rect 20578 5070 20580 5122
rect 20524 5058 20580 5070
rect 20636 5122 20692 5134
rect 20636 5070 20638 5122
rect 20690 5070 20692 5122
rect 20636 4900 20692 5070
rect 20636 4834 20692 4844
rect 20748 4898 20804 4910
rect 20748 4846 20750 4898
rect 20802 4846 20804 4898
rect 19964 4620 20692 4676
rect 19964 4562 20020 4620
rect 19964 4510 19966 4562
rect 20018 4510 20020 4562
rect 19964 4498 20020 4510
rect 19740 4398 19742 4450
rect 19794 4398 19796 4450
rect 19740 4386 19796 4398
rect 20076 4452 20132 4462
rect 20076 4358 20132 4396
rect 20636 4450 20692 4620
rect 20636 4398 20638 4450
rect 20690 4398 20692 4450
rect 20636 4386 20692 4398
rect 18732 4286 18734 4338
rect 18786 4286 18788 4338
rect 18732 4274 18788 4286
rect 20748 4340 20804 4846
rect 21420 4452 21476 4462
rect 21532 4452 21588 6076
rect 21756 6066 21812 6076
rect 21644 5908 21700 5918
rect 21644 5814 21700 5852
rect 22092 5906 22148 5918
rect 22092 5854 22094 5906
rect 22146 5854 22148 5906
rect 21420 4450 21588 4452
rect 21420 4398 21422 4450
rect 21474 4398 21588 4450
rect 21420 4396 21588 4398
rect 21868 5012 21924 5022
rect 21420 4386 21476 4396
rect 20972 4340 21028 4350
rect 20748 4338 21140 4340
rect 20748 4286 20974 4338
rect 21026 4286 21140 4338
rect 20748 4284 21140 4286
rect 20972 4274 21028 4284
rect 14252 4226 14308 4238
rect 14252 4174 14254 4226
rect 14306 4174 14308 4226
rect 14252 4116 14308 4174
rect 13692 4060 14308 4116
rect 19068 4114 19124 4126
rect 19068 4062 19070 4114
rect 19122 4062 19124 4114
rect 13468 3780 13524 3790
rect 13692 3780 13748 4060
rect 13468 3778 13748 3780
rect 13468 3726 13470 3778
rect 13522 3726 13748 3778
rect 13468 3724 13748 3726
rect 19068 3780 19124 4062
rect 20972 4116 21028 4126
rect 20972 4022 21028 4060
rect 13468 3714 13524 3724
rect 19068 3714 19124 3724
rect 13244 3614 13246 3666
rect 13298 3614 13300 3666
rect 13244 3602 13300 3614
rect 13132 3502 13134 3554
rect 13186 3502 13188 3554
rect 4284 3444 4340 3482
rect 4284 3378 4340 3388
rect 6748 3442 6804 3500
rect 13132 3490 13188 3502
rect 21084 3556 21140 4284
rect 21868 4114 21924 4956
rect 22092 4564 22148 5854
rect 22428 5908 22484 5918
rect 22484 5852 22596 5908
rect 22428 5814 22484 5852
rect 22540 5236 22596 5852
rect 22672 5516 22936 5526
rect 22728 5460 22776 5516
rect 22832 5460 22880 5516
rect 22672 5450 22936 5460
rect 22540 5142 22596 5180
rect 23324 5122 23380 6412
rect 23324 5070 23326 5122
rect 23378 5070 23380 5122
rect 23324 5058 23380 5070
rect 23660 5122 23716 6636
rect 24108 6626 24164 6636
rect 24220 6802 24276 12012
rect 25228 11284 25284 11294
rect 24668 10836 24724 10846
rect 24668 10742 24724 10780
rect 24444 9828 24500 9838
rect 24668 9828 24724 9838
rect 24500 9826 24724 9828
rect 24500 9774 24670 9826
rect 24722 9774 24724 9826
rect 24500 9772 24724 9774
rect 24444 9154 24500 9772
rect 24668 9762 24724 9772
rect 24444 9102 24446 9154
rect 24498 9102 24500 9154
rect 24444 9090 24500 9102
rect 24556 9156 24612 9166
rect 24556 8370 24612 9100
rect 24556 8318 24558 8370
rect 24610 8318 24612 8370
rect 24556 7700 24612 8318
rect 25228 9042 25284 11228
rect 25788 11284 25844 11294
rect 26012 11284 26068 14366
rect 26684 14700 26796 14756
rect 26684 13972 26740 14700
rect 26796 14690 26852 14700
rect 26796 14476 26964 14532
rect 26796 14306 26852 14476
rect 26908 14420 26964 14476
rect 27132 14420 27188 15092
rect 28364 14754 28420 14766
rect 28364 14702 28366 14754
rect 28418 14702 28420 14754
rect 28364 14644 28420 14702
rect 28476 14644 28532 14654
rect 28364 14588 28476 14644
rect 28476 14578 28532 14588
rect 27468 14532 27524 14542
rect 27468 14438 27524 14476
rect 28252 14532 28308 14542
rect 28308 14476 28420 14532
rect 28252 14466 28308 14476
rect 26908 14418 27188 14420
rect 26908 14366 27134 14418
rect 27186 14366 27188 14418
rect 26908 14364 27188 14366
rect 26796 14254 26798 14306
rect 26850 14254 26852 14306
rect 26796 14196 26852 14254
rect 26796 14130 26852 14140
rect 26796 13972 26852 13982
rect 26684 13970 26852 13972
rect 26684 13918 26798 13970
rect 26850 13918 26852 13970
rect 26684 13916 26852 13918
rect 26796 13906 26852 13916
rect 27132 13972 27188 14364
rect 28364 14418 28420 14476
rect 28364 14366 28366 14418
rect 28418 14366 28420 14418
rect 27132 13906 27188 13916
rect 27244 14308 27300 14318
rect 27804 14308 27860 14318
rect 27244 14306 27860 14308
rect 27244 14254 27246 14306
rect 27298 14254 27806 14306
rect 27858 14254 27860 14306
rect 27244 14252 27860 14254
rect 26124 13748 26180 13758
rect 26124 12178 26180 13692
rect 26684 13748 26740 13758
rect 26684 13654 26740 13692
rect 26908 13746 26964 13758
rect 26908 13694 26910 13746
rect 26962 13694 26964 13746
rect 26460 13634 26516 13646
rect 26460 13582 26462 13634
rect 26514 13582 26516 13634
rect 26236 13522 26292 13534
rect 26460 13524 26516 13582
rect 26236 13470 26238 13522
rect 26290 13470 26292 13522
rect 26236 12404 26292 13470
rect 26236 12338 26292 12348
rect 26348 13468 26460 13524
rect 26124 12126 26126 12178
rect 26178 12126 26180 12178
rect 26124 12114 26180 12126
rect 26236 11508 26292 11518
rect 26348 11508 26404 13468
rect 26460 13458 26516 13468
rect 26908 13636 26964 13694
rect 26908 12964 26964 13580
rect 27244 13188 27300 14252
rect 27804 14242 27860 14252
rect 27692 13972 27748 13982
rect 27692 13878 27748 13916
rect 27804 13748 27860 13758
rect 27804 13654 27860 13692
rect 27916 13746 27972 13758
rect 27916 13694 27918 13746
rect 27970 13694 27972 13746
rect 27916 13636 27972 13694
rect 28364 13746 28420 14366
rect 28476 14418 28532 14430
rect 28476 14366 28478 14418
rect 28530 14366 28532 14418
rect 28476 13970 28532 14366
rect 28476 13918 28478 13970
rect 28530 13918 28532 13970
rect 28476 13906 28532 13918
rect 28588 13860 28644 15932
rect 29148 13972 29204 18396
rect 29596 18386 29652 18396
rect 29708 17108 29764 18508
rect 30380 17668 30436 20076
rect 30492 20066 30548 20076
rect 30604 20130 30660 20636
rect 30604 20078 30606 20130
rect 30658 20078 30660 20130
rect 30492 19794 30548 19806
rect 30492 19742 30494 19794
rect 30546 19742 30548 19794
rect 30492 18450 30548 19742
rect 30604 19796 30660 20078
rect 30716 20578 30772 20590
rect 30716 20526 30718 20578
rect 30770 20526 30772 20578
rect 30716 20020 30772 20526
rect 30828 20356 30884 22206
rect 31276 22930 31332 22942
rect 31276 22878 31278 22930
rect 31330 22878 31332 22930
rect 31052 21588 31108 21598
rect 31052 21494 31108 21532
rect 31052 20580 31108 20590
rect 31052 20486 31108 20524
rect 30828 20290 30884 20300
rect 30716 19954 30772 19964
rect 30604 19740 30884 19796
rect 30492 18398 30494 18450
rect 30546 18398 30548 18450
rect 30492 18386 30548 18398
rect 30828 18450 30884 19740
rect 31276 19460 31332 22878
rect 31388 21698 31444 22988
rect 31388 21646 31390 21698
rect 31442 21646 31444 21698
rect 31388 21634 31444 21646
rect 31612 20804 31668 25564
rect 32060 25618 32116 25630
rect 32060 25566 32062 25618
rect 32114 25566 32116 25618
rect 32060 25508 32116 25566
rect 32060 25442 32116 25452
rect 31836 25172 31892 25182
rect 31724 25060 31780 25070
rect 31724 24946 31780 25004
rect 31724 24894 31726 24946
rect 31778 24894 31780 24946
rect 31724 24882 31780 24894
rect 31612 20738 31668 20748
rect 31724 23826 31780 23838
rect 31724 23774 31726 23826
rect 31778 23774 31780 23826
rect 31276 19404 31444 19460
rect 31164 19236 31220 19246
rect 31164 19142 31220 19180
rect 30828 18398 30830 18450
rect 30882 18398 30884 18450
rect 30828 18386 30884 18398
rect 30156 17612 30380 17668
rect 29825 17276 30089 17286
rect 29881 17220 29929 17276
rect 29985 17220 30033 17276
rect 29825 17210 30089 17220
rect 29708 17052 30100 17108
rect 29260 16996 29316 17006
rect 29260 16882 29316 16940
rect 29260 16830 29262 16882
rect 29314 16830 29316 16882
rect 29260 16818 29316 16830
rect 29596 16884 29652 16894
rect 29596 16436 29652 16828
rect 29596 16370 29652 16380
rect 30044 16098 30100 17052
rect 30044 16046 30046 16098
rect 30098 16046 30100 16098
rect 30044 16034 30100 16046
rect 30156 15986 30212 17612
rect 30380 17602 30436 17612
rect 30716 18338 30772 18350
rect 30716 18286 30718 18338
rect 30770 18286 30772 18338
rect 30716 16994 30772 18286
rect 31164 18226 31220 18238
rect 31164 18174 31166 18226
rect 31218 18174 31220 18226
rect 31164 17668 31220 18174
rect 31164 17602 31220 17612
rect 30716 16942 30718 16994
rect 30770 16942 30772 16994
rect 30716 16772 30772 16942
rect 31052 16884 31108 16894
rect 30716 16706 30772 16716
rect 30828 16882 31108 16884
rect 30828 16830 31054 16882
rect 31106 16830 31108 16882
rect 30828 16828 31108 16830
rect 30156 15934 30158 15986
rect 30210 15934 30212 15986
rect 30156 15922 30212 15934
rect 30268 16548 30324 16558
rect 29825 15708 30089 15718
rect 29881 15652 29929 15708
rect 29985 15652 30033 15708
rect 29825 15642 30089 15652
rect 30268 15540 30324 16492
rect 30828 16436 30884 16828
rect 31052 16818 31108 16828
rect 31276 16660 31332 16670
rect 30380 16380 30884 16436
rect 31164 16658 31332 16660
rect 31164 16606 31278 16658
rect 31330 16606 31332 16658
rect 31164 16604 31332 16606
rect 30380 16098 30436 16380
rect 31164 16322 31220 16604
rect 31164 16270 31166 16322
rect 31218 16270 31220 16322
rect 31164 16258 31220 16270
rect 30380 16046 30382 16098
rect 30434 16046 30436 16098
rect 30380 16034 30436 16046
rect 30828 15876 30884 15886
rect 30828 15874 31108 15876
rect 30828 15822 30830 15874
rect 30882 15822 31108 15874
rect 30828 15820 31108 15822
rect 30828 15810 30884 15820
rect 29825 14140 30089 14150
rect 29881 14084 29929 14140
rect 29985 14084 30033 14140
rect 29825 14074 30089 14084
rect 29260 13972 29316 13982
rect 28812 13970 29316 13972
rect 28812 13918 29262 13970
rect 29314 13918 29316 13970
rect 28812 13916 29316 13918
rect 28588 13794 28644 13804
rect 28700 13858 28756 13870
rect 28700 13806 28702 13858
rect 28754 13806 28756 13858
rect 28364 13694 28366 13746
rect 28418 13694 28420 13746
rect 28364 13682 28420 13694
rect 27916 13300 27972 13580
rect 28700 13636 28756 13806
rect 28812 13858 28868 13916
rect 29260 13906 29316 13916
rect 28812 13806 28814 13858
rect 28866 13806 28868 13858
rect 28812 13794 28868 13806
rect 30044 13860 30100 13870
rect 30044 13766 30100 13804
rect 30268 13746 30324 15484
rect 30828 15316 30884 15326
rect 30828 15222 30884 15260
rect 31052 15314 31108 15820
rect 31052 15262 31054 15314
rect 31106 15262 31108 15314
rect 31052 15250 31108 15262
rect 30268 13694 30270 13746
rect 30322 13694 30324 13746
rect 30268 13682 30324 13694
rect 30716 14530 30772 14542
rect 30716 14478 30718 14530
rect 30770 14478 30772 14530
rect 30716 13970 30772 14478
rect 30716 13918 30718 13970
rect 30770 13918 30772 13970
rect 28700 13570 28756 13580
rect 29708 13636 29764 13646
rect 29708 13542 29764 13580
rect 26908 12962 27188 12964
rect 26908 12910 26910 12962
rect 26962 12910 27188 12962
rect 26908 12908 27188 12910
rect 26908 12898 26964 12908
rect 26460 12738 26516 12750
rect 26460 12686 26462 12738
rect 26514 12686 26516 12738
rect 26460 12404 26516 12686
rect 26460 12338 26516 12348
rect 26796 11508 26852 11518
rect 26236 11506 27076 11508
rect 26236 11454 26238 11506
rect 26290 11454 26798 11506
rect 26850 11454 27076 11506
rect 26236 11452 27076 11454
rect 26236 11442 26292 11452
rect 26796 11414 26852 11452
rect 25844 11228 26068 11284
rect 26796 11284 26852 11294
rect 25788 11190 25844 11228
rect 26572 11172 26628 11182
rect 25900 11060 25956 11070
rect 25900 10834 25956 11004
rect 25900 10782 25902 10834
rect 25954 10782 25956 10834
rect 25900 10770 25956 10782
rect 26572 10834 26628 11116
rect 26572 10782 26574 10834
rect 26626 10782 26628 10834
rect 26572 10770 26628 10782
rect 25452 10612 25508 10622
rect 25452 10518 25508 10556
rect 26348 10610 26404 10622
rect 26348 10558 26350 10610
rect 26402 10558 26404 10610
rect 26348 10388 26404 10558
rect 26572 10612 26628 10622
rect 26572 10518 26628 10556
rect 26796 10612 26852 11228
rect 26796 10546 26852 10556
rect 26908 10610 26964 10622
rect 26908 10558 26910 10610
rect 26962 10558 26964 10610
rect 26908 10500 26964 10558
rect 26908 10434 26964 10444
rect 26348 9714 26404 10332
rect 26348 9662 26350 9714
rect 26402 9662 26404 9714
rect 26348 9650 26404 9662
rect 27020 10050 27076 11452
rect 27132 11396 27188 12908
rect 27244 12962 27300 13132
rect 27244 12910 27246 12962
rect 27298 12910 27300 12962
rect 27244 12898 27300 12910
rect 27692 13244 27972 13300
rect 27692 12404 27748 13244
rect 28252 13188 28308 13198
rect 28252 13094 28308 13132
rect 29148 13188 29204 13198
rect 28364 13074 28420 13086
rect 28364 13022 28366 13074
rect 28418 13022 28420 13074
rect 27692 12338 27748 12348
rect 28140 12962 28196 12974
rect 28140 12910 28142 12962
rect 28194 12910 28196 12962
rect 28140 12178 28196 12910
rect 28252 12404 28308 12414
rect 28364 12404 28420 13022
rect 28308 12348 28420 12404
rect 29148 12402 29204 13132
rect 30604 12962 30660 12974
rect 30604 12910 30606 12962
rect 30658 12910 30660 12962
rect 30604 12852 30660 12910
rect 30716 12964 30772 13918
rect 31164 14532 31220 14542
rect 30940 13188 30996 13198
rect 30940 13094 30996 13132
rect 30716 12898 30772 12908
rect 31052 12964 31108 12974
rect 31164 12964 31220 14476
rect 31276 13188 31332 16604
rect 31388 16210 31444 19404
rect 31500 17666 31556 17678
rect 31500 17614 31502 17666
rect 31554 17614 31556 17666
rect 31500 16548 31556 17614
rect 31724 17108 31780 23774
rect 31836 21586 31892 25116
rect 32284 24948 32340 25900
rect 32396 25620 32452 25630
rect 32396 25506 32452 25564
rect 32396 25454 32398 25506
rect 32450 25454 32452 25506
rect 32396 25442 32452 25454
rect 32732 25508 32788 25518
rect 32732 25394 32788 25452
rect 32732 25342 32734 25394
rect 32786 25342 32788 25394
rect 32284 24892 32452 24948
rect 32172 24836 32228 24846
rect 32396 24836 32452 24892
rect 32228 24780 32340 24836
rect 32172 24742 32228 24780
rect 32060 24724 32116 24734
rect 31948 24722 32116 24724
rect 31948 24670 32062 24722
rect 32114 24670 32116 24722
rect 31948 24668 32116 24670
rect 31948 23492 32004 24668
rect 32060 24658 32116 24668
rect 32172 24500 32228 24510
rect 31948 23426 32004 23436
rect 32060 24498 32228 24500
rect 32060 24446 32174 24498
rect 32226 24446 32228 24498
rect 32060 24444 32228 24446
rect 32060 23154 32116 24444
rect 32172 24434 32228 24444
rect 32060 23102 32062 23154
rect 32114 23102 32116 23154
rect 32060 23090 32116 23102
rect 31836 21534 31838 21586
rect 31890 21534 31892 21586
rect 31836 21522 31892 21534
rect 32060 22370 32116 22382
rect 32060 22318 32062 22370
rect 32114 22318 32116 22370
rect 31948 21474 32004 21486
rect 31948 21422 31950 21474
rect 32002 21422 32004 21474
rect 31836 20804 31892 20814
rect 31836 20710 31892 20748
rect 31948 18564 32004 21422
rect 32060 19236 32116 22318
rect 32284 21586 32340 24780
rect 32396 24770 32452 24780
rect 32732 23826 32788 25342
rect 32844 25506 32900 25518
rect 32844 25454 32846 25506
rect 32898 25454 32900 25506
rect 32844 25396 32900 25454
rect 32844 23938 32900 25340
rect 33068 24610 33124 26238
rect 33740 26292 33796 26302
rect 33740 26290 33908 26292
rect 33740 26238 33742 26290
rect 33794 26238 33908 26290
rect 33740 26236 33908 26238
rect 33740 26226 33796 26236
rect 33516 26178 33572 26190
rect 33516 26126 33518 26178
rect 33570 26126 33572 26178
rect 33068 24558 33070 24610
rect 33122 24558 33124 24610
rect 33068 24546 33124 24558
rect 33180 24834 33236 24846
rect 33180 24782 33182 24834
rect 33234 24782 33236 24834
rect 33180 24724 33236 24782
rect 33180 24164 33236 24668
rect 33404 24836 33460 24846
rect 33404 24164 33460 24780
rect 33516 24724 33572 26126
rect 33852 25396 33908 26236
rect 34188 26290 34244 26302
rect 34188 26238 34190 26290
rect 34242 26238 34244 26290
rect 34188 26180 34244 26238
rect 35532 26292 35588 26302
rect 33852 25340 34132 25396
rect 33740 25172 33796 25182
rect 33740 24834 33796 25116
rect 34076 24946 34132 25340
rect 34076 24894 34078 24946
rect 34130 24894 34132 24946
rect 34076 24882 34132 24894
rect 33740 24782 33742 24834
rect 33794 24782 33796 24834
rect 33740 24770 33796 24782
rect 33852 24834 33908 24846
rect 33852 24782 33854 24834
rect 33906 24782 33908 24834
rect 33516 24658 33572 24668
rect 33404 24108 33684 24164
rect 33180 24098 33236 24108
rect 33628 24050 33684 24108
rect 33628 23998 33630 24050
rect 33682 23998 33684 24050
rect 33628 23986 33684 23998
rect 32844 23886 32846 23938
rect 32898 23886 32900 23938
rect 32844 23874 32900 23886
rect 32732 23774 32734 23826
rect 32786 23774 32788 23826
rect 32732 23762 32788 23774
rect 33404 23716 33460 23726
rect 32284 21534 32286 21586
rect 32338 21534 32340 21586
rect 32284 21522 32340 21534
rect 32732 22370 32788 22382
rect 32732 22318 32734 22370
rect 32786 22318 32788 22370
rect 32396 21252 32452 21262
rect 32172 20804 32228 20814
rect 32172 20710 32228 20748
rect 32396 20802 32452 21196
rect 32396 20750 32398 20802
rect 32450 20750 32452 20802
rect 32396 20738 32452 20750
rect 32060 19170 32116 19180
rect 32396 19346 32452 19358
rect 32396 19294 32398 19346
rect 32450 19294 32452 19346
rect 31948 18498 32004 18508
rect 32172 17666 32228 17678
rect 32172 17614 32174 17666
rect 32226 17614 32228 17666
rect 31612 17052 31780 17108
rect 32060 17108 32116 17118
rect 31612 16548 31668 17052
rect 32060 16882 32116 17052
rect 32060 16830 32062 16882
rect 32114 16830 32116 16882
rect 32060 16818 32116 16830
rect 32172 16884 32228 17614
rect 32172 16818 32228 16828
rect 31724 16772 31780 16782
rect 31724 16678 31780 16716
rect 31612 16492 31892 16548
rect 31500 16482 31556 16492
rect 31388 16158 31390 16210
rect 31442 16158 31444 16210
rect 31388 15148 31444 16158
rect 31724 15204 31780 15242
rect 31388 15092 31668 15148
rect 31724 15138 31780 15148
rect 31276 13132 31556 13188
rect 31276 12964 31332 12974
rect 31164 12962 31332 12964
rect 31164 12910 31278 12962
rect 31330 12910 31332 12962
rect 31164 12908 31332 12910
rect 30604 12786 30660 12796
rect 29148 12350 29150 12402
rect 29202 12350 29204 12402
rect 28252 12338 28308 12348
rect 29148 12338 29204 12350
rect 29260 12738 29316 12750
rect 29260 12686 29262 12738
rect 29314 12686 29316 12738
rect 28140 12126 28142 12178
rect 28194 12126 28196 12178
rect 27356 12068 27412 12078
rect 27916 12068 27972 12078
rect 27356 12066 27916 12068
rect 27356 12014 27358 12066
rect 27410 12014 27916 12066
rect 27356 12012 27916 12014
rect 27356 12002 27412 12012
rect 27916 11974 27972 12012
rect 27132 11394 27412 11396
rect 27132 11342 27134 11394
rect 27186 11342 27412 11394
rect 27132 11340 27412 11342
rect 27132 11330 27188 11340
rect 27356 10834 27412 11340
rect 27356 10782 27358 10834
rect 27410 10782 27412 10834
rect 27020 9998 27022 10050
rect 27074 9998 27076 10050
rect 27020 9604 27076 9998
rect 26908 9602 27076 9604
rect 26908 9550 27022 9602
rect 27074 9550 27076 9602
rect 26908 9548 27076 9550
rect 25788 9156 25844 9166
rect 25788 9062 25844 9100
rect 26684 9156 26740 9166
rect 26684 9062 26740 9100
rect 25228 8990 25230 9042
rect 25282 8990 25284 9042
rect 25004 8260 25060 8270
rect 25004 8166 25060 8204
rect 25228 8036 25284 8990
rect 25452 9044 25508 9054
rect 26012 9044 26068 9054
rect 25452 8950 25508 8988
rect 25900 9042 26068 9044
rect 25900 8990 26014 9042
rect 26066 8990 26068 9042
rect 25900 8988 26068 8990
rect 25676 8932 25732 8942
rect 25452 8146 25508 8158
rect 25452 8094 25454 8146
rect 25506 8094 25508 8146
rect 25452 8036 25508 8094
rect 24556 7634 24612 7644
rect 24668 7980 25396 8036
rect 24668 7698 24724 7980
rect 24668 7646 24670 7698
rect 24722 7646 24724 7698
rect 24668 7634 24724 7646
rect 25228 7252 25284 7262
rect 25116 7250 25284 7252
rect 25116 7198 25230 7250
rect 25282 7198 25284 7250
rect 25116 7196 25284 7198
rect 24220 6750 24222 6802
rect 24274 6750 24276 6802
rect 23660 5070 23662 5122
rect 23714 5070 23716 5122
rect 23660 5058 23716 5070
rect 23884 6466 23940 6478
rect 23884 6414 23886 6466
rect 23938 6414 23940 6466
rect 23884 5012 23940 6414
rect 23996 5236 24052 5246
rect 24220 5236 24276 6750
rect 23996 5234 24276 5236
rect 23996 5182 23998 5234
rect 24050 5182 24276 5234
rect 23996 5180 24276 5182
rect 24332 6916 24388 6926
rect 23996 5170 24052 5180
rect 23884 4956 24164 5012
rect 22092 4498 22148 4508
rect 22876 4900 22932 4910
rect 22764 4452 22820 4462
rect 22764 4358 22820 4396
rect 22428 4340 22484 4350
rect 21868 4062 21870 4114
rect 21922 4062 21924 4114
rect 21868 4050 21924 4062
rect 22204 4284 22428 4340
rect 21868 3780 21924 3790
rect 21868 3686 21924 3724
rect 22204 3778 22260 4284
rect 22428 4246 22484 4284
rect 22876 4338 22932 4844
rect 23996 4564 24052 4574
rect 23996 4470 24052 4508
rect 24108 4450 24164 4956
rect 24332 4562 24388 6860
rect 25004 6916 25060 6926
rect 25004 6578 25060 6860
rect 25004 6526 25006 6578
rect 25058 6526 25060 6578
rect 25004 6514 25060 6526
rect 25116 6578 25172 7196
rect 25228 7186 25284 7196
rect 25116 6526 25118 6578
rect 25170 6526 25172 6578
rect 24780 6468 24836 6478
rect 24780 6374 24836 6412
rect 24332 4510 24334 4562
rect 24386 4510 24388 4562
rect 24332 4498 24388 4510
rect 24556 4676 24612 4686
rect 24108 4398 24110 4450
rect 24162 4398 24164 4450
rect 22876 4286 22878 4338
rect 22930 4286 22932 4338
rect 22876 4274 22932 4286
rect 23772 4340 23828 4350
rect 23772 4246 23828 4284
rect 23436 4116 23492 4126
rect 23436 4022 23492 4060
rect 23772 4116 23828 4126
rect 23772 4022 23828 4060
rect 24108 4004 24164 4398
rect 22672 3948 22936 3958
rect 22728 3892 22776 3948
rect 22832 3892 22880 3948
rect 24108 3938 24164 3948
rect 22672 3882 22936 3892
rect 22204 3726 22206 3778
rect 22258 3726 22260 3778
rect 22204 3714 22260 3726
rect 23660 3780 23716 3790
rect 23660 3666 23716 3724
rect 23660 3614 23662 3666
rect 23714 3614 23716 3666
rect 23660 3602 23716 3614
rect 21084 3490 21140 3500
rect 21644 3556 21700 3566
rect 21644 3462 21700 3500
rect 24556 3554 24612 4620
rect 24668 4340 24724 4350
rect 25116 4340 25172 6526
rect 25340 6132 25396 7980
rect 25452 7970 25508 7980
rect 25676 7586 25732 8876
rect 25900 8482 25956 8988
rect 26012 8978 26068 8988
rect 26124 9044 26180 9054
rect 26460 9044 26516 9054
rect 25900 8430 25902 8482
rect 25954 8430 25956 8482
rect 25900 8260 25956 8430
rect 25900 8194 25956 8204
rect 26012 8260 26068 8270
rect 26124 8260 26180 8988
rect 26012 8258 26124 8260
rect 26012 8206 26014 8258
rect 26066 8206 26124 8258
rect 26012 8204 26124 8206
rect 26012 8194 26068 8204
rect 26124 8194 26180 8204
rect 26348 9042 26516 9044
rect 26348 8990 26462 9042
rect 26514 8990 26516 9042
rect 26348 8988 26516 8990
rect 25676 7534 25678 7586
rect 25730 7534 25732 7586
rect 25676 7522 25732 7534
rect 25788 8148 25844 8158
rect 25788 7588 25844 8092
rect 25900 8034 25956 8046
rect 25900 7982 25902 8034
rect 25954 7982 25956 8034
rect 25900 7924 25956 7982
rect 25900 7858 25956 7868
rect 26124 8036 26180 8046
rect 25788 7494 25844 7532
rect 26012 7476 26068 7486
rect 26124 7476 26180 7980
rect 26236 7924 26292 7934
rect 26348 7924 26404 8988
rect 26460 8978 26516 8988
rect 26572 8932 26628 8942
rect 26572 8838 26628 8876
rect 26908 8484 26964 9548
rect 27020 9538 27076 9548
rect 27132 10724 27188 10734
rect 27132 9044 27188 10668
rect 27356 10052 27412 10782
rect 28140 11282 28196 12126
rect 28140 11230 28142 11282
rect 28194 11230 28196 11282
rect 28140 10610 28196 11230
rect 28140 10558 28142 10610
rect 28194 10558 28196 10610
rect 28028 10052 28084 10062
rect 28140 10052 28196 10558
rect 27412 9996 27636 10052
rect 27356 9986 27412 9996
rect 27580 9938 27636 9996
rect 27580 9886 27582 9938
rect 27634 9886 27636 9938
rect 27580 9874 27636 9886
rect 28028 10050 28196 10052
rect 28028 9998 28030 10050
rect 28082 9998 28196 10050
rect 28028 9996 28196 9998
rect 28364 12180 28420 12190
rect 28364 10610 28420 12124
rect 29260 12180 29316 12686
rect 30828 12738 30884 12750
rect 30828 12686 30830 12738
rect 30882 12686 30884 12738
rect 29825 12572 30089 12582
rect 29881 12516 29929 12572
rect 29985 12516 30033 12572
rect 29825 12506 30089 12516
rect 29484 12180 29540 12190
rect 29316 12178 29540 12180
rect 29316 12126 29486 12178
rect 29538 12126 29540 12178
rect 29316 12124 29540 12126
rect 29260 12114 29316 12124
rect 29484 12114 29540 12124
rect 29148 11732 29204 11742
rect 28476 11170 28532 11182
rect 28476 11118 28478 11170
rect 28530 11118 28532 11170
rect 28476 10724 28532 11118
rect 28476 10658 28532 10668
rect 28812 11172 28868 11182
rect 28364 10558 28366 10610
rect 28418 10558 28420 10610
rect 28364 10052 28420 10558
rect 28812 10612 28868 11116
rect 29148 10834 29204 11676
rect 30156 11620 30212 11630
rect 30156 11526 30212 11564
rect 30380 11508 30436 11518
rect 30380 11394 30436 11452
rect 30380 11342 30382 11394
rect 30434 11342 30436 11394
rect 30044 11284 30100 11294
rect 30100 11228 30212 11284
rect 29820 11172 29876 11210
rect 30044 11190 30100 11228
rect 29820 11106 29876 11116
rect 29825 11004 30089 11014
rect 29881 10948 29929 11004
rect 29985 10948 30033 11004
rect 29825 10938 30089 10948
rect 29148 10782 29150 10834
rect 29202 10782 29204 10834
rect 29148 10770 29204 10782
rect 29484 10836 29540 10846
rect 29484 10722 29540 10780
rect 29932 10836 29988 10846
rect 29932 10742 29988 10780
rect 29484 10670 29486 10722
rect 29538 10670 29540 10722
rect 29484 10658 29540 10670
rect 30156 10612 30212 11228
rect 30380 10836 30436 11342
rect 30828 11284 30884 12686
rect 31052 12290 31108 12908
rect 31276 12402 31332 12908
rect 31388 12964 31444 12974
rect 31388 12850 31444 12908
rect 31388 12798 31390 12850
rect 31442 12798 31444 12850
rect 31388 12786 31444 12798
rect 31276 12350 31278 12402
rect 31330 12350 31332 12402
rect 31276 12338 31332 12350
rect 31052 12238 31054 12290
rect 31106 12238 31108 12290
rect 31052 12226 31108 12238
rect 31164 12066 31220 12078
rect 31164 12014 31166 12066
rect 31218 12014 31220 12066
rect 31164 11506 31220 12014
rect 31164 11454 31166 11506
rect 31218 11454 31220 11506
rect 31164 11442 31220 11454
rect 31276 11284 31332 11294
rect 30828 11282 31332 11284
rect 30828 11230 31278 11282
rect 31330 11230 31332 11282
rect 30828 11228 31332 11230
rect 31276 11218 31332 11228
rect 30492 10836 30548 10846
rect 30436 10834 30548 10836
rect 30436 10782 30494 10834
rect 30546 10782 30548 10834
rect 30436 10780 30548 10782
rect 30380 10742 30436 10780
rect 30492 10770 30548 10780
rect 31500 10612 31556 13132
rect 30156 10556 30324 10612
rect 28812 10498 28868 10556
rect 28812 10446 28814 10498
rect 28866 10446 28868 10498
rect 28812 10434 28868 10446
rect 28028 9938 28084 9996
rect 28364 9986 28420 9996
rect 29372 10386 29428 10398
rect 29372 10334 29374 10386
rect 29426 10334 29428 10386
rect 28028 9886 28030 9938
rect 28082 9886 28084 9938
rect 28028 9874 28084 9886
rect 27468 9268 27524 9278
rect 27356 9156 27412 9166
rect 27356 9062 27412 9100
rect 26908 8418 26964 8428
rect 27020 8988 27188 9044
rect 26460 8260 26516 8270
rect 26908 8260 26964 8270
rect 26516 8258 26964 8260
rect 26516 8206 26910 8258
rect 26962 8206 26964 8258
rect 26516 8204 26964 8206
rect 26460 8166 26516 8204
rect 26908 8194 26964 8204
rect 26292 7868 26404 7924
rect 26236 7858 26292 7868
rect 26012 7474 26180 7476
rect 26012 7422 26014 7474
rect 26066 7422 26180 7474
rect 26012 7420 26180 7422
rect 26012 7410 26068 7420
rect 26012 6804 26068 6814
rect 25340 6130 25956 6132
rect 25340 6078 25342 6130
rect 25394 6078 25956 6130
rect 25340 6076 25956 6078
rect 25340 6066 25396 6076
rect 25676 5684 25732 5694
rect 25564 5012 25620 5022
rect 25452 5010 25620 5012
rect 25452 4958 25566 5010
rect 25618 4958 25620 5010
rect 25452 4956 25620 4958
rect 25228 4676 25284 4686
rect 25228 4562 25284 4620
rect 25228 4510 25230 4562
rect 25282 4510 25284 4562
rect 25228 4498 25284 4510
rect 25452 4562 25508 4956
rect 25564 4946 25620 4956
rect 25452 4510 25454 4562
rect 25506 4510 25508 4562
rect 24668 4338 25172 4340
rect 24668 4286 24670 4338
rect 24722 4286 25172 4338
rect 24668 4284 25172 4286
rect 24668 4274 24724 4284
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24668 3556 24724 3566
rect 6748 3390 6750 3442
rect 6802 3390 6804 3442
rect 6748 3378 6804 3390
rect 23772 3444 23828 3482
rect 23772 3378 23828 3388
rect 24668 3442 24724 3500
rect 24892 3556 24948 3566
rect 25116 3556 25172 3566
rect 24892 3554 25172 3556
rect 24892 3502 24894 3554
rect 24946 3502 25118 3554
rect 25170 3502 25172 3554
rect 24892 3500 25172 3502
rect 24892 3490 24948 3500
rect 25116 3490 25172 3500
rect 25452 3556 25508 4510
rect 25564 4452 25620 4462
rect 25676 4452 25732 5628
rect 25788 5236 25844 5246
rect 25788 5122 25844 5180
rect 25788 5070 25790 5122
rect 25842 5070 25844 5122
rect 25788 5058 25844 5070
rect 25564 4450 25732 4452
rect 25564 4398 25566 4450
rect 25618 4398 25732 4450
rect 25564 4396 25732 4398
rect 25564 4386 25620 4396
rect 25900 4338 25956 6076
rect 25900 4286 25902 4338
rect 25954 4286 25956 4338
rect 25900 4274 25956 4286
rect 26012 4226 26068 6748
rect 27020 5908 27076 8988
rect 27468 8372 27524 9212
rect 28028 9268 28084 9278
rect 27356 8316 27524 8372
rect 27580 9042 27636 9054
rect 27580 8990 27582 9042
rect 27634 8990 27636 9042
rect 27580 8484 27636 8990
rect 28028 9042 28084 9212
rect 28028 8990 28030 9042
rect 28082 8990 28084 9042
rect 27580 8428 27972 8484
rect 27132 8260 27188 8270
rect 27132 8166 27188 8204
rect 27356 8146 27412 8316
rect 27356 8094 27358 8146
rect 27410 8094 27412 8146
rect 27356 7588 27412 8094
rect 27468 8148 27524 8158
rect 27580 8148 27636 8428
rect 27804 8260 27860 8270
rect 27468 8146 27636 8148
rect 27468 8094 27470 8146
rect 27522 8094 27636 8146
rect 27468 8092 27636 8094
rect 27468 8082 27524 8092
rect 27468 7588 27524 7598
rect 27356 7586 27524 7588
rect 27356 7534 27470 7586
rect 27522 7534 27524 7586
rect 27356 7532 27524 7534
rect 27468 7522 27524 7532
rect 27580 6914 27636 8092
rect 27692 8258 27860 8260
rect 27692 8206 27806 8258
rect 27858 8206 27860 8258
rect 27692 8204 27860 8206
rect 27692 7700 27748 8204
rect 27804 8194 27860 8204
rect 27916 8036 27972 8428
rect 28028 8258 28084 8990
rect 28364 8818 28420 8830
rect 28364 8766 28366 8818
rect 28418 8766 28420 8818
rect 28364 8372 28420 8766
rect 29372 8372 29428 10334
rect 30268 9826 30324 10556
rect 31276 10610 31556 10612
rect 31276 10558 31502 10610
rect 31554 10558 31556 10610
rect 31276 10556 31556 10558
rect 30716 10052 30772 10062
rect 30716 9938 30772 9996
rect 30716 9886 30718 9938
rect 30770 9886 30772 9938
rect 30716 9874 30772 9886
rect 30268 9774 30270 9826
rect 30322 9774 30324 9826
rect 30268 9762 30324 9774
rect 31276 9826 31332 10556
rect 31500 10546 31556 10556
rect 31612 10612 31668 15092
rect 31836 14308 31892 16492
rect 32060 15876 32116 15886
rect 32060 15314 32116 15820
rect 32060 15262 32062 15314
rect 32114 15262 32116 15314
rect 32060 15250 32116 15262
rect 32396 14532 32452 19294
rect 32620 19236 32676 19246
rect 32732 19236 32788 22318
rect 33404 22258 33460 23660
rect 33852 23380 33908 24782
rect 34188 24836 34244 26124
rect 35420 26180 35476 26190
rect 35420 26086 35476 26124
rect 35532 25620 35588 26236
rect 35532 25526 35588 25564
rect 35980 26180 36036 26190
rect 34524 25508 34580 25518
rect 34188 24770 34244 24780
rect 34300 25506 34580 25508
rect 34300 25454 34526 25506
rect 34578 25454 34580 25506
rect 34300 25452 34580 25454
rect 33628 23324 33908 23380
rect 33628 23044 33684 23324
rect 33740 23156 33796 23166
rect 33740 23062 33796 23100
rect 33628 22950 33684 22988
rect 33404 22206 33406 22258
rect 33458 22206 33460 22258
rect 33404 22194 33460 22206
rect 33516 22370 33572 22382
rect 33516 22318 33518 22370
rect 33570 22318 33572 22370
rect 33516 20692 33572 22318
rect 34300 21812 34356 25452
rect 34524 25442 34580 25452
rect 35420 25396 35476 25406
rect 35308 25340 35420 25396
rect 34972 25284 35028 25294
rect 34972 25190 35028 25228
rect 34972 24948 35028 24958
rect 34748 24836 34804 24846
rect 34524 24164 34580 24174
rect 34412 23156 34468 23166
rect 34412 22258 34468 23100
rect 34524 22820 34580 24108
rect 34748 24052 34804 24780
rect 34748 23958 34804 23996
rect 34972 24834 35028 24892
rect 34972 24782 34974 24834
rect 35026 24782 35028 24834
rect 34972 23828 35028 24782
rect 35308 24050 35364 25340
rect 35420 25330 35476 25340
rect 35868 25394 35924 25406
rect 35868 25342 35870 25394
rect 35922 25342 35924 25394
rect 35756 25172 35812 25182
rect 35308 23998 35310 24050
rect 35362 23998 35364 24050
rect 35308 23986 35364 23998
rect 35420 24052 35476 24062
rect 35084 23828 35140 23838
rect 34972 23826 35252 23828
rect 34972 23774 35086 23826
rect 35138 23774 35252 23826
rect 34972 23772 35252 23774
rect 35084 23762 35140 23772
rect 34748 23044 34804 23054
rect 34748 23042 35140 23044
rect 34748 22990 34750 23042
rect 34802 22990 35140 23042
rect 34748 22988 35140 22990
rect 34748 22978 34804 22988
rect 35084 22932 35140 22988
rect 34524 22764 34804 22820
rect 34412 22206 34414 22258
rect 34466 22206 34468 22258
rect 34412 22194 34468 22206
rect 34412 21812 34468 21822
rect 34300 21756 34412 21812
rect 34412 21586 34468 21756
rect 34412 21534 34414 21586
rect 34466 21534 34468 21586
rect 34412 21522 34468 21534
rect 34748 21028 34804 22764
rect 35084 22596 35140 22876
rect 35196 22820 35252 23772
rect 35308 23716 35364 23726
rect 35308 23622 35364 23660
rect 35308 23266 35364 23278
rect 35308 23214 35310 23266
rect 35362 23214 35364 23266
rect 35308 23156 35364 23214
rect 35308 23090 35364 23100
rect 35420 23154 35476 23996
rect 35756 23938 35812 25116
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35756 23874 35812 23886
rect 35868 24946 35924 25342
rect 35868 24894 35870 24946
rect 35922 24894 35924 24946
rect 35868 23940 35924 24894
rect 35980 24050 36036 26124
rect 36092 25506 36148 26348
rect 37436 26402 37492 26414
rect 37436 26350 37438 26402
rect 37490 26350 37492 26402
rect 36204 26292 36260 26302
rect 36204 26198 36260 26236
rect 36316 26068 36372 26078
rect 36092 25454 36094 25506
rect 36146 25454 36148 25506
rect 36092 25442 36148 25454
rect 36204 26066 36372 26068
rect 36204 26014 36318 26066
rect 36370 26014 36372 26066
rect 36204 26012 36372 26014
rect 36204 25508 36260 26012
rect 36316 26002 36372 26012
rect 37436 26068 37492 26350
rect 39116 26404 39172 26414
rect 37436 26002 37492 26012
rect 37996 26290 38052 26302
rect 37996 26238 37998 26290
rect 38050 26238 38052 26290
rect 36979 25900 37243 25910
rect 37035 25844 37083 25900
rect 37139 25844 37187 25900
rect 36979 25834 37243 25844
rect 37548 25730 37604 25742
rect 37548 25678 37550 25730
rect 37602 25678 37604 25730
rect 36092 24164 36148 24174
rect 36204 24164 36260 25452
rect 36428 25508 36484 25518
rect 36428 25414 36484 25452
rect 36988 25506 37044 25518
rect 36988 25454 36990 25506
rect 37042 25454 37044 25506
rect 36316 25284 36372 25294
rect 36316 25190 36372 25228
rect 36988 24948 37044 25454
rect 36988 24882 37044 24892
rect 37212 25506 37268 25518
rect 37212 25454 37214 25506
rect 37266 25454 37268 25506
rect 36092 24162 36260 24164
rect 36092 24110 36094 24162
rect 36146 24110 36260 24162
rect 36092 24108 36260 24110
rect 36428 24836 36484 24846
rect 36428 24722 36484 24780
rect 37212 24836 37268 25454
rect 37548 25508 37604 25678
rect 37212 24770 37268 24780
rect 37436 25172 37492 25182
rect 37436 24834 37492 25116
rect 37436 24782 37438 24834
rect 37490 24782 37492 24834
rect 37436 24770 37492 24782
rect 36428 24670 36430 24722
rect 36482 24670 36484 24722
rect 36092 24098 36148 24108
rect 35980 23998 35982 24050
rect 36034 23998 36036 24050
rect 35980 23986 36036 23998
rect 35868 23874 35924 23884
rect 36428 23716 36484 24670
rect 36979 24332 37243 24342
rect 37035 24276 37083 24332
rect 37139 24276 37187 24332
rect 36979 24266 37243 24276
rect 37548 23826 37604 25452
rect 37996 25172 38052 26238
rect 38556 26180 38612 26190
rect 38556 26178 38948 26180
rect 38556 26126 38558 26178
rect 38610 26126 38948 26178
rect 38556 26124 38948 26126
rect 38556 26114 38612 26124
rect 38780 25508 38836 25518
rect 38892 25508 38948 26124
rect 39004 25508 39060 25518
rect 38892 25506 39060 25508
rect 38892 25454 39006 25506
rect 39058 25454 39060 25506
rect 38892 25452 39060 25454
rect 38780 25284 38836 25452
rect 39004 25442 39060 25452
rect 38668 25228 38836 25284
rect 38668 25172 38724 25228
rect 37996 25106 38052 25116
rect 38556 25116 38724 25172
rect 38556 24722 38612 25116
rect 38556 24670 38558 24722
rect 38610 24670 38612 24722
rect 38556 24658 38612 24670
rect 37884 23940 37940 23950
rect 37884 23938 38164 23940
rect 37884 23886 37886 23938
rect 37938 23886 38164 23938
rect 37884 23884 38164 23886
rect 37884 23874 37940 23884
rect 37548 23774 37550 23826
rect 37602 23774 37604 23826
rect 37548 23762 37604 23774
rect 36428 23650 36484 23660
rect 38108 23604 38164 23884
rect 38108 23538 38164 23548
rect 38556 23714 38612 23726
rect 38556 23662 38558 23714
rect 38610 23662 38612 23714
rect 38220 23266 38276 23278
rect 38220 23214 38222 23266
rect 38274 23214 38276 23266
rect 35420 23102 35422 23154
rect 35474 23102 35476 23154
rect 35196 22764 35364 22820
rect 35196 22596 35252 22606
rect 35084 22594 35252 22596
rect 35084 22542 35198 22594
rect 35250 22542 35252 22594
rect 35084 22540 35252 22542
rect 35196 22530 35252 22540
rect 35308 22372 35364 22764
rect 35196 22316 35364 22372
rect 34860 22258 34916 22270
rect 34860 22206 34862 22258
rect 34914 22206 34916 22258
rect 34860 21252 34916 22206
rect 34916 21196 35140 21252
rect 34860 21186 34916 21196
rect 34860 21028 34916 21038
rect 34748 21026 34916 21028
rect 34748 20974 34862 21026
rect 34914 20974 34916 21026
rect 34748 20972 34916 20974
rect 34860 20962 34916 20972
rect 34524 20914 34580 20926
rect 34524 20862 34526 20914
rect 34578 20862 34580 20914
rect 34524 20804 34580 20862
rect 34524 20738 34580 20748
rect 33516 20626 33572 20636
rect 34188 20692 34244 20702
rect 34188 20598 34244 20636
rect 35084 20692 35140 21196
rect 35084 20598 35140 20636
rect 32620 19234 32788 19236
rect 32620 19182 32622 19234
rect 32674 19182 32788 19234
rect 32620 19180 32788 19182
rect 32844 20578 32900 20590
rect 32844 20526 32846 20578
rect 32898 20526 32900 20578
rect 32620 17890 32676 19180
rect 32620 17838 32622 17890
rect 32674 17838 32676 17890
rect 32620 17826 32676 17838
rect 32508 15314 32564 15326
rect 32508 15262 32510 15314
rect 32562 15262 32564 15314
rect 32508 14980 32564 15262
rect 32844 15148 32900 20526
rect 34412 20578 34468 20590
rect 34972 20580 35028 20590
rect 34412 20526 34414 20578
rect 34466 20526 34468 20578
rect 34188 20356 34244 20366
rect 33068 20020 33124 20030
rect 33068 19926 33124 19964
rect 34188 20018 34244 20300
rect 34188 19966 34190 20018
rect 34242 19966 34244 20018
rect 34188 19954 34244 19966
rect 34412 19460 34468 20526
rect 34412 19394 34468 19404
rect 34636 20578 35028 20580
rect 34636 20526 34974 20578
rect 35026 20526 35028 20578
rect 34636 20524 35028 20526
rect 33516 19236 33572 19246
rect 34076 19236 34132 19246
rect 33180 18450 33236 18462
rect 33180 18398 33182 18450
rect 33234 18398 33236 18450
rect 33068 18226 33124 18238
rect 33068 18174 33070 18226
rect 33122 18174 33124 18226
rect 33068 17220 33124 18174
rect 33068 17154 33124 17164
rect 33180 17668 33236 18398
rect 33404 18452 33460 18462
rect 33404 18358 33460 18396
rect 33292 17668 33348 17678
rect 33180 17666 33348 17668
rect 33180 17614 33294 17666
rect 33346 17614 33348 17666
rect 33180 17612 33348 17614
rect 33068 16996 33124 17006
rect 33180 16996 33236 17612
rect 33292 17602 33348 17612
rect 33516 17108 33572 19180
rect 33964 19234 34132 19236
rect 33964 19182 34078 19234
rect 34130 19182 34132 19234
rect 33964 19180 34132 19182
rect 33852 19124 33908 19134
rect 33852 19030 33908 19068
rect 33852 18452 33908 18462
rect 33964 18452 34020 19180
rect 34076 19170 34132 19180
rect 33852 18450 34020 18452
rect 33852 18398 33854 18450
rect 33906 18398 34020 18450
rect 33852 18396 34020 18398
rect 33516 17042 33572 17052
rect 33628 18226 33684 18238
rect 33628 18174 33630 18226
rect 33682 18174 33684 18226
rect 33124 16940 33236 16996
rect 33068 16902 33124 16940
rect 33292 16884 33348 16894
rect 33628 16884 33684 18174
rect 33348 16828 33684 16884
rect 33740 17220 33796 17230
rect 33292 16790 33348 16828
rect 33516 16660 33572 16670
rect 33516 16566 33572 16604
rect 33740 16658 33796 17164
rect 33740 16606 33742 16658
rect 33794 16606 33796 16658
rect 33740 16212 33796 16606
rect 33852 16660 33908 18396
rect 34524 18338 34580 18350
rect 34524 18286 34526 18338
rect 34578 18286 34580 18338
rect 34524 18116 34580 18286
rect 34524 17556 34580 18060
rect 34524 17490 34580 17500
rect 34300 17108 34356 17118
rect 34636 17108 34692 20524
rect 34972 20514 35028 20524
rect 34972 19460 35028 19470
rect 35028 19404 35140 19460
rect 34972 19394 35028 19404
rect 35084 18674 35140 19404
rect 35196 19458 35252 22316
rect 35308 21812 35364 21822
rect 35308 20018 35364 21756
rect 35420 21700 35476 23102
rect 35756 23156 35812 23166
rect 35420 21634 35476 21644
rect 35532 22146 35588 22158
rect 35532 22094 35534 22146
rect 35586 22094 35588 22146
rect 35308 19966 35310 20018
rect 35362 19966 35364 20018
rect 35308 19954 35364 19966
rect 35308 19796 35364 19806
rect 35364 19740 35476 19796
rect 35308 19730 35364 19740
rect 35196 19406 35198 19458
rect 35250 19406 35252 19458
rect 35196 19394 35252 19406
rect 35084 18622 35086 18674
rect 35138 18622 35140 18674
rect 35084 18610 35140 18622
rect 34300 16994 34356 17052
rect 34300 16942 34302 16994
rect 34354 16942 34356 16994
rect 34300 16930 34356 16942
rect 34412 17052 34692 17108
rect 34748 18564 34804 18574
rect 33852 16594 33908 16604
rect 33740 16146 33796 16156
rect 34188 15540 34244 15550
rect 33964 15316 34020 15326
rect 33964 15222 34020 15260
rect 34188 15314 34244 15484
rect 34188 15262 34190 15314
rect 34242 15262 34244 15314
rect 34188 15250 34244 15262
rect 34412 15316 34468 17052
rect 34636 16884 34692 16894
rect 34636 16790 34692 16828
rect 34748 15540 34804 18508
rect 34972 18562 35028 18574
rect 34972 18510 34974 18562
rect 35026 18510 35028 18562
rect 34972 18340 35028 18510
rect 35196 18452 35252 18462
rect 35252 18396 35364 18452
rect 35196 18386 35252 18396
rect 34860 18284 35028 18340
rect 35084 18340 35140 18350
rect 34860 18116 34916 18284
rect 35084 18228 35140 18284
rect 35196 18228 35252 18238
rect 34860 18050 34916 18060
rect 34972 18226 35252 18228
rect 34972 18174 35198 18226
rect 35250 18174 35252 18226
rect 34972 18172 35252 18174
rect 34972 17108 35028 18172
rect 35196 18162 35252 18172
rect 34972 16882 35028 17052
rect 35196 16996 35252 17006
rect 35308 16996 35364 18396
rect 35196 16994 35364 16996
rect 35196 16942 35198 16994
rect 35250 16942 35364 16994
rect 35196 16940 35364 16942
rect 35196 16930 35252 16940
rect 34972 16830 34974 16882
rect 35026 16830 35028 16882
rect 34972 16818 35028 16830
rect 35084 16770 35140 16782
rect 35084 16718 35086 16770
rect 35138 16718 35140 16770
rect 34860 16212 34916 16222
rect 35084 16212 35140 16718
rect 35084 16156 35252 16212
rect 34860 15986 34916 16156
rect 34860 15934 34862 15986
rect 34914 15934 34916 15986
rect 34860 15922 34916 15934
rect 35084 15988 35140 15998
rect 35084 15894 35140 15932
rect 34972 15874 35028 15886
rect 34972 15822 34974 15874
rect 35026 15822 35028 15874
rect 34748 15484 34916 15540
rect 34636 15316 34692 15326
rect 34860 15316 34916 15484
rect 34412 15314 34580 15316
rect 34412 15262 34414 15314
rect 34466 15262 34580 15314
rect 34412 15260 34580 15262
rect 34412 15250 34468 15260
rect 33516 15202 33572 15214
rect 33516 15150 33518 15202
rect 33570 15150 33572 15202
rect 32844 15092 33124 15148
rect 32508 14914 32564 14924
rect 33068 14642 33124 15092
rect 33516 14980 33572 15150
rect 34524 15148 34580 15260
rect 34636 15314 34916 15316
rect 34636 15262 34638 15314
rect 34690 15262 34916 15314
rect 34636 15260 34916 15262
rect 34636 15250 34692 15260
rect 34524 15092 34804 15148
rect 33516 14914 33572 14924
rect 33068 14590 33070 14642
rect 33122 14590 33124 14642
rect 32396 14466 32452 14476
rect 32956 14530 33012 14542
rect 32956 14478 32958 14530
rect 33010 14478 33012 14530
rect 32956 14308 33012 14478
rect 31836 14252 33012 14308
rect 32956 12852 33012 14252
rect 33068 13188 33124 14590
rect 33068 12964 33124 13132
rect 33516 14754 33572 14766
rect 33516 14702 33518 14754
rect 33570 14702 33572 14754
rect 33292 12964 33348 12974
rect 33068 12962 33348 12964
rect 33068 12910 33294 12962
rect 33346 12910 33348 12962
rect 33068 12908 33348 12910
rect 33292 12898 33348 12908
rect 32956 12786 33012 12796
rect 32060 12628 32116 12638
rect 32060 11620 32116 12572
rect 32060 11554 32116 11564
rect 32956 12292 33012 12302
rect 32956 11284 33012 12236
rect 33516 12180 33572 14702
rect 34748 14642 34804 15092
rect 34748 14590 34750 14642
rect 34802 14590 34804 14642
rect 34748 14578 34804 14590
rect 34860 14530 34916 15260
rect 34972 15316 35028 15822
rect 34972 15222 35028 15260
rect 35196 15540 35252 16156
rect 35196 15314 35252 15484
rect 35196 15262 35198 15314
rect 35250 15262 35252 15314
rect 35196 15250 35252 15262
rect 34860 14478 34862 14530
rect 34914 14478 34916 14530
rect 34860 14466 34916 14478
rect 34412 14420 34468 14430
rect 34412 13970 34468 14364
rect 34748 14308 34804 14318
rect 34748 14306 34916 14308
rect 34748 14254 34750 14306
rect 34802 14254 34916 14306
rect 34748 14252 34916 14254
rect 34748 14242 34804 14252
rect 34412 13918 34414 13970
rect 34466 13918 34468 13970
rect 34412 13906 34468 13918
rect 34748 13636 34804 13646
rect 34860 13636 34916 14252
rect 34972 13636 35028 13646
rect 34860 13634 35028 13636
rect 34860 13582 34974 13634
rect 35026 13582 35028 13634
rect 34860 13580 35028 13582
rect 34748 13542 34804 13580
rect 34972 13524 35028 13580
rect 34972 13458 35028 13468
rect 35308 12962 35364 12974
rect 35308 12910 35310 12962
rect 35362 12910 35364 12962
rect 33852 12852 33908 12862
rect 33852 12758 33908 12796
rect 35084 12852 35140 12862
rect 34972 12740 35028 12750
rect 34972 12646 35028 12684
rect 34972 12404 35028 12414
rect 34860 12348 34972 12404
rect 33516 12114 33572 12124
rect 34188 12180 34244 12190
rect 34188 12086 34244 12124
rect 32284 11282 33012 11284
rect 32284 11230 32958 11282
rect 33010 11230 33012 11282
rect 32284 11228 33012 11230
rect 32284 10722 32340 11228
rect 32956 11218 33012 11228
rect 33180 11282 33236 11294
rect 33180 11230 33182 11282
rect 33234 11230 33236 11282
rect 33180 11060 33236 11230
rect 33180 10994 33236 11004
rect 32284 10670 32286 10722
rect 32338 10670 32340 10722
rect 32284 10658 32340 10670
rect 31724 10612 31780 10622
rect 31612 10610 31780 10612
rect 31612 10558 31726 10610
rect 31778 10558 31780 10610
rect 31612 10556 31780 10558
rect 31276 9774 31278 9826
rect 31330 9774 31332 9826
rect 31276 9762 31332 9774
rect 31612 9826 31668 10556
rect 31724 10546 31780 10556
rect 34860 10610 34916 12348
rect 34972 12338 35028 12348
rect 35084 12292 35140 12796
rect 35084 12198 35140 12236
rect 35308 12180 35364 12910
rect 35308 12114 35364 12124
rect 35420 12068 35476 19740
rect 35532 17444 35588 22094
rect 35756 19908 35812 23100
rect 36876 23156 36932 23194
rect 36876 23090 36932 23100
rect 37100 23156 37156 23166
rect 37100 23154 37380 23156
rect 37100 23102 37102 23154
rect 37154 23102 37380 23154
rect 37100 23100 37380 23102
rect 37100 23090 37156 23100
rect 36316 23044 36372 23054
rect 36316 22950 36372 22988
rect 35980 22932 36036 22942
rect 35868 22876 35980 22932
rect 35868 21586 35924 22876
rect 35980 22838 36036 22876
rect 37212 22932 37268 22970
rect 37212 22866 37268 22876
rect 36979 22764 37243 22774
rect 37035 22708 37083 22764
rect 37139 22708 37187 22764
rect 36979 22698 37243 22708
rect 36204 22596 36260 22606
rect 36260 22540 36372 22596
rect 36204 22530 36260 22540
rect 35868 21534 35870 21586
rect 35922 21534 35924 21586
rect 35868 21522 35924 21534
rect 36092 20692 36148 20702
rect 36092 20018 36148 20636
rect 36316 20468 36372 22540
rect 36988 22260 37044 22270
rect 36428 21700 36484 21710
rect 36428 21028 36484 21644
rect 36988 21698 37044 22204
rect 36988 21646 36990 21698
rect 37042 21646 37044 21698
rect 36988 21634 37044 21646
rect 37324 21588 37380 23100
rect 37660 23044 37716 23054
rect 37660 22950 37716 22988
rect 38108 23044 38164 23054
rect 38108 22482 38164 22988
rect 38108 22430 38110 22482
rect 38162 22430 38164 22482
rect 38108 22418 38164 22430
rect 37324 21522 37380 21532
rect 37548 22372 37604 22382
rect 37548 21586 37604 22316
rect 38220 22372 38276 23214
rect 38556 22820 38612 23662
rect 39116 23604 39172 26348
rect 40124 26404 40180 26414
rect 40124 26310 40180 26348
rect 41356 26290 41412 26302
rect 41356 26238 41358 26290
rect 41410 26238 41412 26290
rect 39900 26180 39956 26190
rect 39900 26086 39956 26124
rect 40236 26180 40292 26190
rect 40236 25060 40292 26124
rect 41356 25396 41412 26238
rect 48636 26290 48692 26302
rect 48636 26238 48638 26290
rect 48690 26238 48692 26290
rect 46844 26180 46900 26190
rect 46844 26086 46900 26124
rect 47628 26178 47684 26190
rect 47628 26126 47630 26178
rect 47682 26126 47684 26178
rect 42700 26068 42756 26078
rect 42700 26066 43092 26068
rect 42700 26014 42702 26066
rect 42754 26014 43092 26066
rect 42700 26012 43092 26014
rect 42700 26002 42756 26012
rect 42140 25618 42196 25630
rect 42140 25566 42142 25618
rect 42194 25566 42196 25618
rect 41356 25330 41412 25340
rect 41804 25506 41860 25518
rect 41804 25454 41806 25506
rect 41858 25454 41860 25506
rect 40236 24994 40292 25004
rect 39676 24946 39732 24958
rect 41804 24948 41860 25454
rect 39676 24894 39678 24946
rect 39730 24894 39732 24946
rect 39564 24724 39620 24734
rect 39564 24630 39620 24668
rect 39340 24610 39396 24622
rect 39340 24558 39342 24610
rect 39394 24558 39396 24610
rect 39228 23940 39284 23950
rect 39228 23846 39284 23884
rect 38556 22754 38612 22764
rect 39004 22930 39060 22942
rect 39004 22878 39006 22930
rect 39058 22878 39060 22930
rect 39004 22372 39060 22878
rect 38220 22278 38276 22316
rect 38780 22316 39004 22372
rect 38556 22148 38612 22158
rect 37548 21534 37550 21586
rect 37602 21534 37604 21586
rect 36428 20914 36484 20972
rect 36428 20862 36430 20914
rect 36482 20862 36484 20914
rect 36428 20850 36484 20862
rect 36764 21362 36820 21374
rect 36764 21310 36766 21362
rect 36818 21310 36820 21362
rect 36316 20412 36484 20468
rect 36316 20244 36372 20254
rect 36316 20130 36372 20188
rect 36316 20078 36318 20130
rect 36370 20078 36372 20130
rect 36316 20066 36372 20078
rect 36092 19966 36094 20018
rect 36146 19966 36148 20018
rect 36092 19954 36148 19966
rect 36204 20020 36260 20030
rect 35756 19842 35812 19852
rect 35644 19796 35700 19806
rect 35644 19702 35700 19740
rect 36092 19460 36148 19470
rect 35868 19236 35924 19246
rect 35868 19142 35924 19180
rect 36092 19122 36148 19404
rect 36204 19458 36260 19964
rect 36204 19406 36206 19458
rect 36258 19406 36260 19458
rect 36204 19394 36260 19406
rect 36092 19070 36094 19122
rect 36146 19070 36148 19122
rect 36092 19058 36148 19070
rect 35868 18788 35924 18798
rect 35868 18674 35924 18732
rect 35868 18622 35870 18674
rect 35922 18622 35924 18674
rect 35756 18562 35812 18574
rect 35756 18510 35758 18562
rect 35810 18510 35812 18562
rect 35756 18452 35812 18510
rect 35756 18386 35812 18396
rect 35868 18340 35924 18622
rect 36092 18452 36148 18462
rect 36092 18358 36148 18396
rect 36316 18450 36372 18462
rect 36316 18398 36318 18450
rect 36370 18398 36372 18450
rect 35924 18284 36036 18340
rect 35868 18274 35924 18284
rect 35980 17780 36036 18284
rect 35980 17724 36260 17780
rect 35532 17378 35588 17388
rect 35756 17556 35812 17566
rect 35756 17106 35812 17500
rect 35756 17054 35758 17106
rect 35810 17054 35812 17106
rect 35756 17042 35812 17054
rect 36204 16994 36260 17724
rect 36316 17220 36372 18398
rect 36316 17154 36372 17164
rect 36204 16942 36206 16994
rect 36258 16942 36260 16994
rect 36204 16930 36260 16942
rect 36092 16882 36148 16894
rect 36092 16830 36094 16882
rect 36146 16830 36148 16882
rect 36092 15988 36148 16830
rect 36428 16212 36484 20412
rect 36652 19124 36708 19134
rect 36652 18450 36708 19068
rect 36652 18398 36654 18450
rect 36706 18398 36708 18450
rect 36652 18386 36708 18398
rect 36540 18340 36596 18350
rect 36540 18246 36596 18284
rect 36764 16996 36820 21310
rect 36979 21196 37243 21206
rect 37035 21140 37083 21196
rect 37139 21140 37187 21196
rect 36979 21130 37243 21140
rect 36988 21028 37044 21038
rect 36988 20690 37044 20972
rect 36988 20638 36990 20690
rect 37042 20638 37044 20690
rect 36988 20626 37044 20638
rect 37212 20802 37268 20814
rect 37212 20750 37214 20802
rect 37266 20750 37268 20802
rect 37212 20244 37268 20750
rect 37212 20178 37268 20188
rect 37324 19906 37380 19918
rect 37324 19854 37326 19906
rect 37378 19854 37380 19906
rect 36979 19628 37243 19638
rect 37035 19572 37083 19628
rect 37139 19572 37187 19628
rect 36979 19562 37243 19572
rect 37100 19234 37156 19246
rect 37100 19182 37102 19234
rect 37154 19182 37156 19234
rect 37100 18788 37156 19182
rect 37100 18722 37156 18732
rect 37212 19124 37268 19134
rect 37100 18562 37156 18574
rect 37100 18510 37102 18562
rect 37154 18510 37156 18562
rect 37100 18452 37156 18510
rect 37100 18386 37156 18396
rect 37212 18450 37268 19068
rect 37212 18398 37214 18450
rect 37266 18398 37268 18450
rect 37212 18386 37268 18398
rect 36979 18060 37243 18070
rect 37035 18004 37083 18060
rect 37139 18004 37187 18060
rect 36979 17994 37243 18004
rect 36652 16940 36820 16996
rect 37100 17556 37156 17566
rect 36652 16324 36708 16940
rect 37100 16882 37156 17500
rect 37100 16830 37102 16882
rect 37154 16830 37156 16882
rect 37100 16818 37156 16830
rect 36764 16770 36820 16782
rect 36764 16718 36766 16770
rect 36818 16718 36820 16770
rect 36764 16660 36820 16718
rect 36764 16594 36820 16604
rect 36979 16492 37243 16502
rect 37035 16436 37083 16492
rect 37139 16436 37187 16492
rect 36979 16426 37243 16436
rect 36652 16268 37044 16324
rect 36428 16118 36484 16156
rect 36988 16100 37044 16268
rect 36988 16006 37044 16044
rect 36092 15922 36148 15932
rect 37100 15538 37156 15550
rect 37100 15486 37102 15538
rect 37154 15486 37156 15538
rect 36988 15314 37044 15326
rect 36988 15262 36990 15314
rect 37042 15262 37044 15314
rect 36988 15204 37044 15262
rect 36988 15138 37044 15148
rect 35644 15090 35700 15102
rect 35644 15038 35646 15090
rect 35698 15038 35700 15090
rect 35644 13972 35700 15038
rect 35868 15092 35924 15102
rect 35756 14980 35812 14990
rect 35756 14530 35812 14924
rect 35756 14478 35758 14530
rect 35810 14478 35812 14530
rect 35756 14466 35812 14478
rect 35868 14420 35924 15036
rect 37100 15092 37156 15486
rect 37100 15026 37156 15036
rect 37324 15316 37380 19854
rect 37548 19346 37604 21534
rect 38332 21588 38388 21598
rect 38332 21494 38388 21532
rect 38556 20914 38612 22092
rect 38780 21586 38836 22316
rect 39004 22306 39060 22316
rect 38780 21534 38782 21586
rect 38834 21534 38836 21586
rect 38780 21522 38836 21534
rect 38556 20862 38558 20914
rect 38610 20862 38612 20914
rect 38556 20850 38612 20862
rect 38780 20804 38836 20814
rect 38780 20710 38836 20748
rect 38892 20132 38948 20142
rect 37884 20020 37940 20030
rect 37884 19926 37940 19964
rect 38892 19908 38948 20076
rect 38892 19814 38948 19852
rect 37548 19294 37550 19346
rect 37602 19294 37604 19346
rect 37548 19282 37604 19294
rect 37772 19796 37828 19806
rect 37548 17668 37604 17678
rect 37548 17574 37604 17612
rect 37772 17666 37828 19740
rect 39004 19234 39060 19246
rect 39004 19182 39006 19234
rect 39058 19182 39060 19234
rect 38780 18452 38836 18462
rect 38780 18358 38836 18396
rect 39004 17780 39060 19182
rect 39004 17714 39060 17724
rect 39116 17778 39172 23548
rect 39340 23828 39396 24558
rect 39340 23156 39396 23772
rect 39228 23100 39396 23156
rect 39676 23380 39732 24894
rect 41692 24892 41860 24948
rect 41692 24724 41748 24892
rect 41020 23938 41076 23950
rect 41020 23886 41022 23938
rect 41074 23886 41076 23938
rect 41020 23828 41076 23886
rect 41020 23762 41076 23772
rect 41692 23826 41748 24668
rect 41692 23774 41694 23826
rect 41746 23774 41748 23826
rect 41692 23762 41748 23774
rect 42028 24722 42084 24734
rect 42028 24670 42030 24722
rect 42082 24670 42084 24722
rect 39228 18674 39284 23100
rect 39676 22484 39732 23324
rect 40572 23604 40628 23614
rect 40348 23156 40404 23166
rect 39900 23044 39956 23054
rect 39900 22950 39956 22988
rect 39676 22418 39732 22428
rect 40348 22482 40404 23100
rect 40348 22430 40350 22482
rect 40402 22430 40404 22482
rect 40348 22418 40404 22430
rect 40012 22372 40068 22382
rect 40012 22278 40068 22316
rect 40236 21474 40292 21486
rect 40236 21422 40238 21474
rect 40290 21422 40292 21474
rect 40236 21364 40292 21422
rect 40236 21298 40292 21308
rect 40348 20690 40404 20702
rect 40348 20638 40350 20690
rect 40402 20638 40404 20690
rect 39340 20020 39396 20030
rect 39676 20020 39732 20030
rect 39340 19906 39396 19964
rect 39340 19854 39342 19906
rect 39394 19854 39396 19906
rect 39340 19124 39396 19854
rect 39340 19058 39396 19068
rect 39564 20018 39732 20020
rect 39564 19966 39678 20018
rect 39730 19966 39732 20018
rect 39564 19964 39732 19966
rect 39228 18622 39230 18674
rect 39282 18622 39284 18674
rect 39228 18610 39284 18622
rect 39564 17892 39620 19964
rect 39676 19954 39732 19964
rect 40236 20020 40292 20030
rect 40236 19926 40292 19964
rect 40348 19908 40404 20638
rect 40236 19124 40292 19134
rect 39564 17826 39620 17836
rect 39676 18676 39732 18686
rect 39116 17726 39118 17778
rect 39170 17726 39172 17778
rect 39116 17714 39172 17726
rect 37772 17614 37774 17666
rect 37826 17614 37828 17666
rect 37772 17602 37828 17614
rect 37548 17444 37604 17454
rect 37548 16994 37604 17388
rect 37548 16942 37550 16994
rect 37602 16942 37604 16994
rect 37548 16100 37604 16942
rect 38892 16882 38948 16894
rect 38892 16830 38894 16882
rect 38946 16830 38948 16882
rect 37772 16660 37828 16670
rect 37772 16210 37828 16604
rect 37772 16158 37774 16210
rect 37826 16158 37828 16210
rect 37772 16146 37828 16158
rect 38108 16658 38164 16670
rect 38108 16606 38110 16658
rect 38162 16606 38164 16658
rect 38108 16212 38164 16606
rect 38108 16156 38500 16212
rect 37660 16100 37716 16110
rect 37548 16098 37716 16100
rect 37548 16046 37662 16098
rect 37714 16046 37716 16098
rect 37548 16044 37716 16046
rect 37660 16034 37716 16044
rect 37884 16100 37940 16110
rect 36979 14924 37243 14934
rect 37035 14868 37083 14924
rect 37139 14868 37187 14924
rect 36979 14858 37243 14868
rect 35868 14326 35924 14364
rect 36988 14532 37044 14542
rect 36092 14308 36148 14318
rect 35980 14306 36148 14308
rect 35980 14254 36094 14306
rect 36146 14254 36148 14306
rect 35980 14252 36148 14254
rect 35644 13916 35924 13972
rect 35756 13746 35812 13758
rect 35756 13694 35758 13746
rect 35810 13694 35812 13746
rect 35756 13524 35812 13694
rect 35868 13636 35924 13916
rect 35868 13542 35924 13580
rect 35756 13458 35812 13468
rect 35868 12962 35924 12974
rect 35868 12910 35870 12962
rect 35922 12910 35924 12962
rect 35756 12852 35812 12862
rect 35756 12758 35812 12796
rect 35420 12002 35476 12012
rect 35532 12738 35588 12750
rect 35532 12686 35534 12738
rect 35586 12686 35588 12738
rect 35532 11844 35588 12686
rect 35868 12740 35924 12910
rect 35868 12178 35924 12684
rect 35980 12404 36036 14252
rect 36092 14242 36148 14252
rect 36204 14308 36260 14318
rect 36092 13860 36148 13870
rect 36092 13766 36148 13804
rect 35980 12338 36036 12348
rect 35868 12126 35870 12178
rect 35922 12126 35924 12178
rect 35868 12114 35924 12126
rect 34860 10558 34862 10610
rect 34914 10558 34916 10610
rect 33740 9940 33796 9950
rect 31612 9774 31614 9826
rect 31666 9774 31668 9826
rect 31612 9762 31668 9774
rect 33628 9884 33740 9940
rect 32844 9716 32900 9726
rect 32844 9622 32900 9660
rect 30604 9602 30660 9614
rect 30604 9550 30606 9602
rect 30658 9550 30660 9602
rect 29825 9436 30089 9446
rect 29881 9380 29929 9436
rect 29985 9380 30033 9436
rect 29825 9370 30089 9380
rect 29372 8316 29540 8372
rect 28364 8306 28420 8316
rect 28028 8206 28030 8258
rect 28082 8206 28084 8258
rect 28028 8194 28084 8206
rect 28140 8146 28196 8158
rect 28140 8094 28142 8146
rect 28194 8094 28196 8146
rect 28140 8036 28196 8094
rect 28588 8148 28644 8158
rect 29148 8148 29204 8158
rect 28588 8146 29204 8148
rect 28588 8094 28590 8146
rect 28642 8094 29150 8146
rect 29202 8094 29204 8146
rect 28588 8092 29204 8094
rect 28588 8082 28644 8092
rect 29148 8082 29204 8092
rect 29372 8148 29428 8158
rect 29372 8054 29428 8092
rect 27916 7980 28196 8036
rect 27692 7474 27748 7644
rect 28252 7476 28308 7486
rect 27692 7422 27694 7474
rect 27746 7422 27748 7474
rect 27692 7410 27748 7422
rect 28140 7420 28252 7476
rect 27916 7364 27972 7374
rect 27916 6916 27972 7308
rect 27580 6862 27582 6914
rect 27634 6862 27636 6914
rect 27580 6850 27636 6862
rect 27692 6914 27972 6916
rect 27692 6862 27918 6914
rect 27970 6862 27972 6914
rect 27692 6860 27972 6862
rect 27692 6132 27748 6860
rect 27916 6850 27972 6860
rect 28140 6802 28196 7420
rect 28252 7382 28308 7420
rect 28924 7476 28980 7486
rect 28924 7382 28980 7420
rect 28140 6750 28142 6802
rect 28194 6750 28196 6802
rect 28140 6738 28196 6750
rect 29036 7250 29092 7262
rect 29036 7198 29038 7250
rect 29090 7198 29092 7250
rect 28252 6132 28308 6142
rect 28812 6132 28868 6142
rect 27356 6076 28196 6132
rect 27356 6018 27412 6076
rect 27356 5966 27358 6018
rect 27410 5966 27412 6018
rect 27356 5954 27412 5966
rect 27020 5842 27076 5852
rect 27020 5684 27076 5694
rect 27020 5590 27076 5628
rect 27244 5236 27300 5246
rect 27244 5142 27300 5180
rect 27132 4900 27188 4910
rect 27132 4806 27188 4844
rect 27356 4898 27412 4910
rect 27356 4846 27358 4898
rect 27410 4846 27412 4898
rect 26684 4452 26740 4462
rect 26684 4358 26740 4396
rect 27132 4340 27188 4350
rect 27356 4340 27412 4846
rect 26012 4174 26014 4226
rect 26066 4174 26068 4226
rect 26012 4162 26068 4174
rect 26796 4338 27412 4340
rect 26796 4286 27134 4338
rect 27186 4286 27412 4338
rect 26796 4284 27412 4286
rect 27468 4900 27524 4910
rect 26796 4226 26852 4284
rect 27132 4274 27188 4284
rect 26796 4174 26798 4226
rect 26850 4174 26852 4226
rect 26796 4162 26852 4174
rect 26460 4116 26516 4126
rect 26460 4022 26516 4060
rect 27356 4116 27412 4126
rect 27468 4116 27524 4844
rect 27692 4562 27748 6076
rect 27804 5908 27860 5918
rect 27804 5814 27860 5852
rect 28140 5348 28196 6076
rect 28308 6076 28420 6132
rect 28252 6038 28308 6076
rect 28252 5348 28308 5358
rect 28140 5346 28308 5348
rect 28140 5294 28254 5346
rect 28306 5294 28308 5346
rect 28140 5292 28308 5294
rect 28252 5282 28308 5292
rect 27804 5122 27860 5134
rect 27804 5070 27806 5122
rect 27858 5070 27860 5122
rect 27804 4900 27860 5070
rect 28140 5124 28196 5134
rect 28364 5124 28420 6076
rect 28812 6038 28868 6076
rect 29036 5460 29092 7198
rect 29484 6916 29540 8316
rect 29708 8260 29764 8270
rect 29708 8166 29764 8204
rect 29596 8034 29652 8046
rect 29596 7982 29598 8034
rect 29650 7982 29652 8034
rect 29596 7028 29652 7982
rect 29825 7868 30089 7878
rect 29881 7812 29929 7868
rect 29985 7812 30033 7868
rect 29825 7802 30089 7812
rect 29932 7476 29988 7486
rect 29932 7382 29988 7420
rect 30268 7476 30324 7486
rect 30268 7382 30324 7420
rect 29596 6972 29876 7028
rect 29484 6860 29764 6916
rect 29036 5394 29092 5404
rect 29596 6580 29652 6590
rect 29596 6132 29652 6524
rect 28476 5348 28532 5358
rect 28476 5254 28532 5292
rect 29596 5346 29652 6076
rect 29596 5294 29598 5346
rect 29650 5294 29652 5346
rect 29596 5282 29652 5294
rect 29708 5348 29764 6860
rect 29820 6692 29876 6972
rect 30604 6804 30660 9550
rect 30828 9602 30884 9614
rect 30828 9550 30830 9602
rect 30882 9550 30884 9602
rect 30828 8932 30884 9550
rect 31052 8932 31108 8942
rect 30828 8930 31220 8932
rect 30828 8878 31054 8930
rect 31106 8878 31220 8930
rect 30828 8876 31220 8878
rect 31052 8866 31108 8876
rect 31164 8484 31220 8876
rect 31276 8484 31332 8494
rect 31164 8428 31276 8484
rect 31276 8418 31332 8428
rect 31052 8372 31108 8382
rect 31052 8258 31108 8316
rect 31836 8372 31892 8382
rect 31836 8278 31892 8316
rect 33404 8372 33460 8382
rect 31052 8206 31054 8258
rect 31106 8206 31108 8258
rect 31052 8194 31108 8206
rect 31164 8260 31220 8270
rect 31164 8146 31220 8204
rect 32732 8260 32788 8270
rect 32732 8166 32788 8204
rect 33404 8258 33460 8316
rect 33516 8372 33572 8382
rect 33628 8372 33684 9884
rect 33740 9874 33796 9884
rect 34300 9828 34356 9838
rect 34860 9828 34916 10558
rect 34300 9826 34916 9828
rect 34300 9774 34302 9826
rect 34354 9774 34916 9826
rect 34300 9772 34916 9774
rect 34972 11788 35588 11844
rect 34972 10722 35028 11788
rect 34972 10670 34974 10722
rect 35026 10670 35028 10722
rect 34300 9762 34356 9772
rect 34188 9714 34244 9726
rect 34188 9662 34190 9714
rect 34242 9662 34244 9714
rect 34188 9604 34244 9662
rect 34972 9604 35028 10670
rect 35196 11172 35252 11182
rect 36204 11172 36260 14252
rect 36764 13748 36820 13758
rect 36988 13748 37044 14476
rect 36764 13746 37044 13748
rect 36764 13694 36766 13746
rect 36818 13694 37044 13746
rect 36764 13692 37044 13694
rect 36428 12740 36484 12750
rect 35196 9826 35252 11116
rect 35196 9774 35198 9826
rect 35250 9774 35252 9826
rect 35196 9762 35252 9774
rect 35868 11116 36260 11172
rect 36316 11172 36372 11182
rect 34188 9548 35028 9604
rect 35196 8820 35252 8830
rect 35084 8764 35196 8820
rect 35084 8482 35140 8764
rect 35196 8754 35252 8764
rect 35084 8430 35086 8482
rect 35138 8430 35140 8482
rect 35084 8418 35140 8430
rect 33516 8370 33684 8372
rect 33516 8318 33518 8370
rect 33570 8318 33684 8370
rect 33516 8316 33684 8318
rect 33516 8306 33572 8316
rect 33404 8206 33406 8258
rect 33458 8206 33460 8258
rect 33404 8194 33460 8206
rect 34076 8258 34132 8270
rect 34076 8206 34078 8258
rect 34130 8206 34132 8258
rect 31164 8094 31166 8146
rect 31218 8094 31220 8146
rect 30828 7588 30884 7598
rect 31164 7588 31220 8094
rect 31612 8146 31668 8158
rect 31612 8094 31614 8146
rect 31666 8094 31668 8146
rect 31388 8036 31444 8046
rect 31388 8034 31556 8036
rect 31388 7982 31390 8034
rect 31442 7982 31556 8034
rect 31388 7980 31556 7982
rect 31388 7970 31444 7980
rect 30828 7586 31220 7588
rect 30828 7534 30830 7586
rect 30882 7534 31220 7586
rect 30828 7532 31220 7534
rect 30828 7522 30884 7532
rect 30604 6738 30660 6748
rect 30828 6916 30884 6926
rect 29820 6626 29876 6636
rect 29825 6300 30089 6310
rect 29881 6244 29929 6300
rect 29985 6244 30033 6300
rect 29825 6234 30089 6244
rect 28140 5122 28420 5124
rect 28140 5070 28142 5122
rect 28194 5070 28420 5122
rect 28140 5068 28420 5070
rect 29708 5122 29764 5292
rect 30604 5460 30660 5470
rect 30604 5234 30660 5404
rect 30604 5182 30606 5234
rect 30658 5182 30660 5234
rect 30604 5170 30660 5182
rect 29708 5070 29710 5122
rect 29762 5070 29764 5122
rect 28140 5058 28196 5068
rect 29708 5058 29764 5070
rect 30828 5122 30884 6860
rect 31500 6804 31556 7980
rect 31612 7028 31668 8094
rect 32508 8148 32564 8158
rect 32508 8054 32564 8092
rect 33292 8148 33348 8158
rect 32172 8034 32228 8046
rect 32172 7982 32174 8034
rect 32226 7982 32228 8034
rect 32172 7476 32228 7982
rect 33068 8036 33124 8046
rect 33068 7942 33124 7980
rect 32172 7410 32228 7420
rect 31612 6962 31668 6972
rect 33068 7252 33124 7262
rect 31500 6748 31780 6804
rect 31724 5906 31780 6748
rect 31724 5854 31726 5906
rect 31778 5854 31780 5906
rect 31724 5842 31780 5854
rect 31948 6692 32004 6702
rect 31948 5906 32004 6636
rect 33068 6690 33124 7196
rect 33068 6638 33070 6690
rect 33122 6638 33124 6690
rect 33068 6626 33124 6638
rect 32732 6580 32788 6590
rect 32508 6578 32788 6580
rect 32508 6526 32734 6578
rect 32786 6526 32788 6578
rect 32508 6524 32788 6526
rect 32396 6468 32452 6478
rect 31948 5854 31950 5906
rect 32002 5854 32004 5906
rect 31948 5842 32004 5854
rect 32284 6412 32396 6468
rect 31500 5684 31556 5694
rect 30828 5070 30830 5122
rect 30882 5070 30884 5122
rect 29148 5012 29204 5022
rect 28924 5010 29204 5012
rect 28924 4958 29150 5010
rect 29202 4958 29204 5010
rect 28924 4956 29204 4958
rect 28140 4900 28196 4910
rect 27804 4898 28196 4900
rect 27804 4846 28142 4898
rect 28194 4846 28196 4898
rect 27804 4844 28196 4846
rect 28140 4834 28196 4844
rect 27692 4510 27694 4562
rect 27746 4510 27748 4562
rect 27692 4498 27748 4510
rect 28476 4564 28532 4574
rect 28700 4564 28756 4574
rect 28476 4562 28700 4564
rect 28476 4510 28478 4562
rect 28530 4510 28700 4562
rect 28476 4508 28700 4510
rect 28476 4498 28532 4508
rect 28700 4498 28756 4508
rect 28364 4338 28420 4350
rect 28364 4286 28366 4338
rect 28418 4286 28420 4338
rect 28364 4228 28420 4286
rect 28588 4340 28644 4350
rect 28588 4246 28644 4284
rect 28364 4162 28420 4172
rect 28924 4228 28980 4956
rect 29148 4946 29204 4956
rect 29372 5010 29428 5022
rect 30828 5012 30884 5070
rect 29372 4958 29374 5010
rect 29426 4958 29428 5010
rect 29260 4898 29316 4910
rect 29260 4846 29262 4898
rect 29314 4846 29316 4898
rect 29260 4676 29316 4846
rect 29036 4620 29316 4676
rect 29036 4338 29092 4620
rect 29372 4452 29428 4958
rect 30604 4956 30884 5012
rect 30940 5460 30996 5470
rect 29825 4732 30089 4742
rect 29881 4676 29929 4732
rect 29985 4676 30033 4732
rect 29825 4666 30089 4676
rect 29372 4386 29428 4396
rect 30604 4450 30660 4956
rect 30604 4398 30606 4450
rect 30658 4398 30660 4450
rect 30604 4386 30660 4398
rect 29036 4286 29038 4338
rect 29090 4286 29092 4338
rect 29036 4274 29092 4286
rect 30828 4340 30884 4350
rect 30940 4340 30996 5404
rect 31500 5234 31556 5628
rect 32172 5684 32228 5694
rect 32172 5590 32228 5628
rect 31500 5182 31502 5234
rect 31554 5182 31556 5234
rect 31500 5170 31556 5182
rect 32172 5124 32228 5134
rect 32284 5124 32340 6412
rect 32396 6374 32452 6412
rect 32228 5068 32340 5124
rect 32396 5908 32452 5918
rect 32508 5908 32564 6524
rect 32732 6514 32788 6524
rect 32844 6468 32900 6478
rect 32844 6374 32900 6412
rect 32396 5906 32564 5908
rect 32396 5854 32398 5906
rect 32450 5854 32564 5906
rect 32396 5852 32564 5854
rect 33292 6018 33348 8092
rect 33628 8148 33684 8158
rect 33628 8054 33684 8092
rect 34076 8148 34132 8206
rect 35868 8258 35924 11116
rect 36316 10722 36372 11116
rect 36316 10670 36318 10722
rect 36370 10670 36372 10722
rect 36316 10658 36372 10670
rect 36428 9940 36484 12684
rect 36764 12402 36820 13692
rect 36979 13356 37243 13366
rect 37035 13300 37083 13356
rect 37139 13300 37187 13356
rect 36979 13290 37243 13300
rect 37324 12962 37380 15260
rect 37884 15314 37940 16044
rect 38108 15426 38164 16156
rect 38108 15374 38110 15426
rect 38162 15374 38164 15426
rect 38108 15362 38164 15374
rect 38220 15986 38276 15998
rect 38220 15934 38222 15986
rect 38274 15934 38276 15986
rect 37884 15262 37886 15314
rect 37938 15262 37940 15314
rect 37884 15250 37940 15262
rect 37884 14642 37940 14654
rect 37884 14590 37886 14642
rect 37938 14590 37940 14642
rect 37884 14532 37940 14590
rect 37884 14466 37940 14476
rect 37996 14530 38052 14542
rect 37996 14478 37998 14530
rect 38050 14478 38052 14530
rect 37548 14196 37604 14206
rect 37996 14196 38052 14478
rect 37436 14140 37548 14196
rect 37436 13746 37492 14140
rect 37548 14130 37604 14140
rect 37884 14140 38052 14196
rect 38220 14530 38276 15934
rect 38220 14478 38222 14530
rect 38274 14478 38276 14530
rect 38220 14196 38276 14478
rect 38332 15202 38388 15214
rect 38332 15150 38334 15202
rect 38386 15150 38388 15202
rect 38332 14420 38388 15150
rect 38332 14354 38388 14364
rect 37436 13694 37438 13746
rect 37490 13694 37492 13746
rect 37436 13682 37492 13694
rect 37884 13860 37940 14140
rect 38220 14130 38276 14140
rect 37884 13634 37940 13804
rect 37884 13582 37886 13634
rect 37938 13582 37940 13634
rect 37884 13570 37940 13582
rect 37996 13636 38052 13646
rect 37324 12910 37326 12962
rect 37378 12910 37380 12962
rect 37324 12898 37380 12910
rect 37436 13524 37492 13534
rect 36764 12350 36766 12402
rect 36818 12350 36820 12402
rect 36764 12338 36820 12350
rect 37436 12290 37492 13468
rect 37548 12962 37604 12974
rect 37548 12910 37550 12962
rect 37602 12910 37604 12962
rect 37548 12852 37604 12910
rect 37772 12964 37828 12974
rect 37772 12870 37828 12908
rect 37660 12852 37716 12862
rect 37548 12850 37716 12852
rect 37548 12798 37662 12850
rect 37714 12798 37716 12850
rect 37548 12796 37716 12798
rect 37660 12516 37716 12796
rect 37660 12450 37716 12460
rect 37436 12238 37438 12290
rect 37490 12238 37492 12290
rect 37436 12226 37492 12238
rect 37996 12178 38052 13580
rect 38444 13636 38500 16156
rect 38780 16100 38836 16110
rect 38892 16100 38948 16830
rect 39676 16884 39732 18620
rect 39788 17668 39844 17678
rect 40236 17668 40292 19068
rect 40348 18340 40404 19852
rect 40572 19346 40628 23548
rect 41244 23156 41300 23166
rect 41244 23062 41300 23100
rect 41580 23154 41636 23166
rect 41580 23102 41582 23154
rect 41634 23102 41636 23154
rect 41356 23042 41412 23054
rect 41356 22990 41358 23042
rect 41410 22990 41412 23042
rect 41020 22820 41076 22830
rect 41020 22370 41076 22764
rect 41020 22318 41022 22370
rect 41074 22318 41076 22370
rect 41020 22306 41076 22318
rect 41356 22148 41412 22990
rect 41468 22484 41524 22494
rect 41468 22390 41524 22428
rect 41356 22082 41412 22092
rect 41580 21700 41636 23102
rect 42028 23156 42084 24670
rect 42140 23828 42196 25566
rect 42700 25396 42756 25406
rect 42700 25302 42756 25340
rect 42364 24722 42420 24734
rect 42364 24670 42366 24722
rect 42418 24670 42420 24722
rect 42252 24612 42308 24622
rect 42252 24518 42308 24556
rect 42140 23762 42196 23772
rect 42028 23090 42084 23100
rect 42252 23156 42308 23166
rect 42252 23062 42308 23100
rect 42364 22148 42420 24670
rect 42700 24724 42756 24734
rect 42700 24630 42756 24668
rect 43036 24722 43092 26012
rect 47628 25732 47684 26126
rect 48076 26180 48132 26190
rect 48076 26086 48132 26124
rect 48636 26180 48692 26238
rect 47684 25676 47908 25732
rect 47628 25666 47684 25676
rect 47516 25620 47572 25630
rect 45388 25508 45444 25518
rect 45276 25506 45444 25508
rect 45276 25454 45390 25506
rect 45442 25454 45444 25506
rect 45276 25452 45444 25454
rect 44492 25396 44548 25406
rect 43036 24670 43038 24722
rect 43090 24670 43092 24722
rect 42924 24612 42980 24622
rect 42924 24518 42980 24556
rect 42924 24052 42980 24062
rect 43036 24052 43092 24670
rect 42924 24050 43092 24052
rect 42924 23998 42926 24050
rect 42978 23998 43092 24050
rect 42924 23996 43092 23998
rect 42924 23986 42980 23996
rect 42812 23938 42868 23950
rect 42812 23886 42814 23938
rect 42866 23886 42868 23938
rect 42812 23156 42868 23886
rect 42924 23156 42980 23166
rect 42812 23100 42924 23156
rect 42924 23062 42980 23100
rect 43036 23042 43092 23996
rect 43260 25282 43316 25294
rect 43260 25230 43262 25282
rect 43314 25230 43316 25282
rect 43260 24722 43316 25230
rect 44132 25116 44396 25126
rect 44188 25060 44236 25116
rect 44292 25060 44340 25116
rect 44132 25050 44396 25060
rect 43260 24670 43262 24722
rect 43314 24670 43316 24722
rect 43260 24612 43316 24670
rect 43260 23604 43316 24556
rect 44492 24610 44548 25340
rect 45164 25394 45220 25406
rect 45164 25342 45166 25394
rect 45218 25342 45220 25394
rect 44716 25284 44772 25294
rect 44716 24834 44772 25228
rect 45164 25284 45220 25342
rect 45276 25396 45332 25452
rect 45388 25442 45444 25452
rect 46508 25506 46564 25518
rect 46508 25454 46510 25506
rect 46562 25454 46564 25506
rect 45276 25330 45332 25340
rect 45164 25218 45220 25228
rect 44716 24782 44718 24834
rect 44770 24782 44772 24834
rect 44716 24770 44772 24782
rect 45948 24724 46004 24734
rect 45948 24630 46004 24668
rect 46508 24724 46564 25454
rect 47516 24724 47572 25564
rect 47852 25396 47908 25676
rect 48636 25506 48692 26124
rect 48636 25454 48638 25506
rect 48690 25454 48692 25506
rect 48636 25442 48692 25454
rect 47852 24946 47908 25340
rect 48188 25284 48244 25294
rect 48188 25190 48244 25228
rect 48972 25284 49028 25294
rect 47852 24894 47854 24946
rect 47906 24894 47908 24946
rect 47852 24882 47908 24894
rect 47516 24668 47684 24724
rect 46508 24658 46564 24668
rect 44492 24558 44494 24610
rect 44546 24558 44548 24610
rect 44492 24546 44548 24558
rect 47292 24500 47348 24510
rect 47516 24500 47572 24510
rect 47292 24498 47572 24500
rect 47292 24446 47294 24498
rect 47346 24446 47518 24498
rect 47570 24446 47572 24498
rect 47292 24444 47572 24446
rect 47292 24434 47348 24444
rect 47516 24434 47572 24444
rect 46844 23940 46900 23950
rect 46844 23846 46900 23884
rect 47180 23938 47236 23950
rect 47180 23886 47182 23938
rect 47234 23886 47236 23938
rect 44268 23828 44324 23838
rect 44492 23828 44548 23838
rect 44268 23826 44492 23828
rect 44268 23774 44270 23826
rect 44322 23774 44492 23826
rect 44268 23772 44492 23774
rect 44268 23762 44324 23772
rect 43260 23538 43316 23548
rect 44132 23548 44396 23558
rect 44188 23492 44236 23548
rect 44292 23492 44340 23548
rect 44132 23482 44396 23492
rect 43036 22990 43038 23042
rect 43090 22990 43092 23042
rect 43036 22978 43092 22990
rect 43596 23044 43652 23054
rect 43596 22370 43652 22988
rect 44268 22484 44324 22494
rect 43596 22318 43598 22370
rect 43650 22318 43652 22370
rect 42364 22082 42420 22092
rect 42924 22148 42980 22158
rect 42980 22092 43092 22148
rect 42924 22082 42980 22092
rect 40572 19294 40574 19346
rect 40626 19294 40628 19346
rect 40460 19122 40516 19134
rect 40460 19070 40462 19122
rect 40514 19070 40516 19122
rect 40460 18676 40516 19070
rect 40460 18610 40516 18620
rect 40348 18246 40404 18284
rect 39788 17666 40292 17668
rect 39788 17614 39790 17666
rect 39842 17614 40292 17666
rect 39788 17612 40292 17614
rect 39788 17602 39844 17612
rect 40236 17106 40292 17612
rect 40236 17054 40238 17106
rect 40290 17054 40292 17106
rect 40236 17042 40292 17054
rect 40348 17780 40404 17790
rect 40124 16884 40180 16894
rect 39676 16882 40180 16884
rect 39676 16830 40126 16882
rect 40178 16830 40180 16882
rect 39676 16828 40180 16830
rect 39228 16772 39284 16782
rect 38836 16044 39060 16100
rect 38780 16006 38836 16044
rect 39004 15538 39060 16044
rect 39228 15986 39284 16716
rect 39228 15934 39230 15986
rect 39282 15934 39284 15986
rect 39228 15922 39284 15934
rect 39452 16770 39508 16782
rect 39452 16718 39454 16770
rect 39506 16718 39508 16770
rect 39004 15486 39006 15538
rect 39058 15486 39060 15538
rect 39004 15474 39060 15486
rect 39340 15204 39396 15242
rect 39340 15138 39396 15148
rect 38668 14754 38724 14766
rect 38668 14702 38670 14754
rect 38722 14702 38724 14754
rect 38668 14196 38724 14702
rect 39452 14532 39508 16718
rect 40124 15876 40180 16828
rect 40348 16212 40404 17724
rect 40460 17108 40516 17118
rect 40460 17014 40516 17052
rect 40460 16212 40516 16222
rect 40348 16210 40516 16212
rect 40348 16158 40462 16210
rect 40514 16158 40516 16210
rect 40348 16156 40516 16158
rect 40236 15876 40292 15886
rect 40124 15874 40292 15876
rect 40124 15822 40238 15874
rect 40290 15822 40292 15874
rect 40124 15820 40292 15822
rect 40236 15540 40292 15820
rect 40236 15474 40292 15484
rect 40348 15316 40404 16156
rect 40460 16146 40516 16156
rect 40012 15260 40404 15316
rect 40012 15204 40068 15260
rect 40572 15148 40628 19294
rect 40796 21644 41636 21700
rect 42140 21700 42196 21710
rect 42140 21698 42308 21700
rect 42140 21646 42142 21698
rect 42194 21646 42308 21698
rect 42140 21644 42308 21646
rect 40796 17556 40852 21644
rect 42140 21634 42196 21644
rect 42028 21586 42084 21598
rect 42028 21534 42030 21586
rect 42082 21534 42084 21586
rect 41132 21474 41188 21486
rect 41132 21422 41134 21474
rect 41186 21422 41188 21474
rect 41132 20804 41188 21422
rect 41468 21474 41524 21486
rect 41468 21422 41470 21474
rect 41522 21422 41524 21474
rect 41468 20916 41524 21422
rect 42028 21364 42084 21534
rect 41468 20860 41972 20916
rect 41020 20802 41188 20804
rect 41020 20750 41134 20802
rect 41186 20750 41188 20802
rect 41020 20748 41188 20750
rect 40908 17780 40964 17790
rect 41020 17780 41076 20748
rect 41132 20738 41188 20748
rect 41916 20802 41972 20860
rect 41916 20750 41918 20802
rect 41970 20750 41972 20802
rect 41804 20692 41860 20702
rect 41468 19908 41524 19918
rect 41468 19906 41636 19908
rect 41468 19854 41470 19906
rect 41522 19854 41636 19906
rect 41468 19852 41636 19854
rect 41468 19842 41524 19852
rect 41132 19234 41188 19246
rect 41132 19182 41134 19234
rect 41186 19182 41188 19234
rect 41132 19124 41188 19182
rect 41132 19058 41188 19068
rect 41468 18676 41524 18686
rect 41468 18582 41524 18620
rect 41244 18564 41300 18574
rect 41244 18470 41300 18508
rect 41356 18338 41412 18350
rect 41356 18286 41358 18338
rect 41410 18286 41412 18338
rect 41244 18116 41300 18126
rect 40908 17778 41020 17780
rect 40908 17726 40910 17778
rect 40962 17726 41020 17778
rect 40908 17724 41020 17726
rect 40908 17714 40964 17724
rect 41020 17686 41076 17724
rect 41132 18060 41244 18116
rect 40796 17500 41076 17556
rect 41020 17106 41076 17500
rect 41020 17054 41022 17106
rect 41074 17054 41076 17106
rect 41020 16548 41076 17054
rect 41132 16882 41188 18060
rect 41244 18050 41300 18060
rect 41356 17668 41412 18286
rect 41580 18340 41636 19852
rect 41692 19236 41748 19246
rect 41692 18674 41748 19180
rect 41804 19234 41860 20636
rect 41804 19182 41806 19234
rect 41858 19182 41860 19234
rect 41804 19170 41860 19182
rect 41692 18622 41694 18674
rect 41746 18622 41748 18674
rect 41692 18610 41748 18622
rect 41916 19124 41972 20750
rect 42028 20804 42084 21308
rect 42140 21028 42196 21038
rect 42140 20934 42196 20972
rect 42028 20738 42084 20748
rect 42252 20244 42308 21644
rect 42364 21586 42420 21598
rect 42364 21534 42366 21586
rect 42418 21534 42420 21586
rect 42364 20580 42420 21534
rect 42364 20514 42420 20524
rect 42700 20802 42756 20814
rect 42700 20750 42702 20802
rect 42754 20750 42756 20802
rect 42364 20244 42420 20254
rect 42252 20188 42364 20244
rect 42364 20178 42420 20188
rect 42028 20020 42084 20030
rect 42028 19926 42084 19964
rect 42364 20020 42420 20030
rect 42700 20020 42756 20750
rect 42364 20018 42756 20020
rect 42364 19966 42366 20018
rect 42418 19966 42756 20018
rect 42364 19964 42756 19966
rect 42812 20802 42868 20814
rect 42812 20750 42814 20802
rect 42866 20750 42868 20802
rect 42812 20020 42868 20750
rect 42364 19796 42420 19964
rect 42812 19954 42868 19964
rect 42364 19730 42420 19740
rect 42924 19908 42980 19918
rect 41916 18564 41972 19068
rect 42924 18676 42980 19852
rect 43036 19122 43092 22092
rect 43596 21588 43652 22318
rect 43372 21532 43596 21588
rect 43260 19908 43316 19918
rect 43260 19814 43316 19852
rect 43148 19236 43204 19246
rect 43372 19236 43428 21532
rect 43596 21522 43652 21532
rect 43932 22428 44268 22484
rect 43708 21474 43764 21486
rect 43708 21422 43710 21474
rect 43762 21422 43764 21474
rect 43708 21028 43764 21422
rect 43708 20962 43764 20972
rect 43820 20244 43876 20254
rect 43820 20130 43876 20188
rect 43820 20078 43822 20130
rect 43874 20078 43876 20130
rect 43820 20066 43876 20078
rect 43932 20132 43988 22428
rect 44268 22390 44324 22428
rect 44044 22258 44100 22270
rect 44044 22206 44046 22258
rect 44098 22206 44100 22258
rect 44044 22148 44100 22206
rect 44492 22260 44548 23772
rect 47068 23826 47124 23838
rect 47068 23774 47070 23826
rect 47122 23774 47124 23826
rect 46284 23714 46340 23726
rect 46284 23662 46286 23714
rect 46338 23662 46340 23714
rect 44604 23042 44660 23054
rect 44604 22990 44606 23042
rect 44658 22990 44660 23042
rect 44604 22372 44660 22990
rect 44828 22372 44884 22382
rect 44604 22316 44828 22372
rect 44492 22204 44772 22260
rect 44044 22082 44100 22092
rect 44132 21980 44396 21990
rect 44188 21924 44236 21980
rect 44292 21924 44340 21980
rect 44132 21914 44396 21924
rect 44044 21586 44100 21598
rect 44044 21534 44046 21586
rect 44098 21534 44100 21586
rect 44044 21476 44100 21534
rect 44716 21586 44772 22204
rect 44716 21534 44718 21586
rect 44770 21534 44772 21586
rect 44716 21522 44772 21534
rect 44044 21410 44100 21420
rect 44492 20804 44548 20814
rect 44044 20692 44100 20702
rect 44044 20598 44100 20636
rect 44132 20412 44396 20422
rect 44188 20356 44236 20412
rect 44292 20356 44340 20412
rect 44132 20346 44396 20356
rect 44380 20244 44436 20254
rect 44156 20132 44212 20142
rect 43932 20130 44212 20132
rect 43932 20078 44158 20130
rect 44210 20078 44212 20130
rect 43932 20076 44212 20078
rect 43148 19234 43428 19236
rect 43148 19182 43150 19234
rect 43202 19182 43428 19234
rect 43148 19180 43428 19182
rect 43932 19460 43988 19470
rect 43148 19170 43204 19180
rect 43036 19070 43038 19122
rect 43090 19070 43092 19122
rect 43036 19058 43092 19070
rect 42812 18620 42980 18676
rect 42812 18564 42868 18620
rect 41916 18508 42532 18564
rect 41804 18340 41860 18350
rect 41580 18284 41804 18340
rect 41580 18116 41636 18284
rect 41804 18274 41860 18284
rect 42140 18338 42196 18350
rect 42140 18286 42142 18338
rect 42194 18286 42196 18338
rect 42140 18228 42196 18286
rect 42140 18162 42196 18172
rect 42252 18228 42308 18238
rect 42252 18226 42420 18228
rect 42252 18174 42254 18226
rect 42306 18174 42420 18226
rect 42252 18172 42420 18174
rect 42252 18162 42308 18172
rect 41580 18050 41636 18060
rect 42252 17892 42308 17902
rect 42252 17798 42308 17836
rect 41692 17780 41748 17790
rect 41468 17668 41524 17678
rect 41356 17666 41524 17668
rect 41356 17614 41470 17666
rect 41522 17614 41524 17666
rect 41356 17612 41524 17614
rect 41468 17602 41524 17612
rect 41692 17666 41748 17724
rect 41692 17614 41694 17666
rect 41746 17614 41748 17666
rect 41692 17602 41748 17614
rect 41804 17778 41860 17790
rect 41804 17726 41806 17778
rect 41858 17726 41860 17778
rect 41132 16830 41134 16882
rect 41186 16830 41188 16882
rect 41132 16818 41188 16830
rect 41244 17554 41300 17566
rect 41244 17502 41246 17554
rect 41298 17502 41300 17554
rect 41244 17108 41300 17502
rect 41804 17444 41860 17726
rect 41916 17668 41972 17678
rect 41916 17666 42308 17668
rect 41916 17614 41918 17666
rect 41970 17614 42308 17666
rect 41916 17612 42308 17614
rect 41916 17602 41972 17612
rect 41244 16770 41300 17052
rect 41580 17388 41860 17444
rect 42252 17444 42308 17612
rect 41580 16884 41636 17388
rect 42140 17108 42196 17118
rect 41580 16818 41636 16828
rect 42028 17052 42140 17108
rect 42028 16772 42084 17052
rect 42140 17014 42196 17052
rect 42252 16996 42308 17388
rect 42364 17108 42420 18172
rect 42476 17442 42532 18508
rect 42812 18450 42868 18508
rect 42812 18398 42814 18450
rect 42866 18398 42868 18450
rect 42812 17892 42868 18398
rect 42924 18452 42980 18462
rect 43596 18452 43652 18462
rect 43932 18452 43988 19404
rect 44156 19236 44212 20076
rect 44156 19170 44212 19180
rect 44380 19012 44436 20188
rect 44492 20018 44548 20748
rect 44492 19966 44494 20018
rect 44546 19966 44548 20018
rect 44492 19954 44548 19966
rect 44380 18956 44548 19012
rect 44132 18844 44396 18854
rect 44188 18788 44236 18844
rect 44292 18788 44340 18844
rect 44132 18778 44396 18788
rect 42924 18358 42980 18396
rect 43036 18450 43988 18452
rect 43036 18398 43598 18450
rect 43650 18398 43988 18450
rect 43036 18396 43988 18398
rect 42812 17826 42868 17836
rect 42476 17390 42478 17442
rect 42530 17390 42532 17442
rect 42476 17332 42532 17390
rect 42476 17266 42532 17276
rect 42588 17778 42644 17790
rect 42588 17726 42590 17778
rect 42642 17726 42644 17778
rect 42588 17220 42644 17726
rect 43036 17554 43092 18396
rect 43596 18386 43652 18396
rect 43260 18116 43316 18126
rect 43260 17890 43316 18060
rect 43260 17838 43262 17890
rect 43314 17838 43316 17890
rect 43260 17826 43316 17838
rect 43036 17502 43038 17554
rect 43090 17502 43092 17554
rect 43036 17490 43092 17502
rect 43148 17444 43204 17454
rect 43148 17350 43204 17388
rect 42588 17164 43652 17220
rect 42364 17052 43540 17108
rect 42252 16940 42532 16996
rect 42476 16882 42532 16940
rect 42476 16830 42478 16882
rect 42530 16830 42532 16882
rect 42476 16818 42532 16830
rect 42588 16884 42644 16894
rect 41244 16718 41246 16770
rect 41298 16718 41300 16770
rect 41244 16706 41300 16718
rect 41692 16716 42084 16772
rect 41020 16492 41524 16548
rect 41132 15484 41412 15540
rect 40908 15316 40964 15326
rect 41132 15316 41188 15484
rect 40964 15314 41188 15316
rect 40964 15262 41134 15314
rect 41186 15262 41188 15314
rect 40964 15260 41188 15262
rect 40908 15250 40964 15260
rect 41132 15250 41188 15260
rect 41244 15316 41300 15326
rect 39564 14644 39620 14654
rect 39564 14550 39620 14588
rect 39340 14476 39508 14532
rect 39228 14420 39284 14430
rect 39228 14326 39284 14364
rect 38444 13570 38500 13580
rect 38556 14140 38668 14196
rect 38556 12962 38612 14140
rect 38668 14102 38724 14140
rect 38556 12910 38558 12962
rect 38610 12910 38612 12962
rect 38556 12898 38612 12910
rect 39228 13524 39284 13534
rect 37996 12126 37998 12178
rect 38050 12126 38052 12178
rect 37996 12114 38052 12126
rect 38668 12516 38724 12526
rect 38332 12068 38388 12078
rect 36979 11788 37243 11798
rect 36764 11732 36820 11742
rect 37035 11732 37083 11788
rect 37139 11732 37187 11788
rect 36979 11722 37243 11732
rect 36764 11508 36820 11676
rect 36764 11442 36820 11452
rect 38220 11172 38276 11182
rect 38220 11078 38276 11116
rect 37772 10836 37828 10846
rect 37660 10388 37716 10398
rect 37660 10294 37716 10332
rect 36979 10220 37243 10230
rect 37035 10164 37083 10220
rect 37139 10164 37187 10220
rect 36979 10154 37243 10164
rect 37772 10052 37828 10780
rect 38332 10836 38388 12012
rect 38668 11396 38724 12460
rect 39004 11396 39060 11406
rect 39228 11396 39284 13468
rect 38668 11394 38948 11396
rect 38668 11342 38670 11394
rect 38722 11342 38948 11394
rect 38668 11340 38948 11342
rect 38668 11330 38724 11340
rect 38892 11172 38948 11340
rect 39004 11394 39284 11396
rect 39004 11342 39006 11394
rect 39058 11342 39284 11394
rect 39004 11340 39284 11342
rect 39004 11330 39060 11340
rect 38892 11116 39172 11172
rect 38332 10742 38388 10780
rect 39116 10610 39172 11116
rect 39228 10724 39284 11340
rect 39340 11284 39396 14476
rect 39900 14420 39956 14430
rect 39452 14306 39508 14318
rect 39452 14254 39454 14306
rect 39506 14254 39508 14306
rect 39452 14196 39508 14254
rect 39452 14130 39508 14140
rect 39564 13860 39620 13870
rect 39564 13634 39620 13804
rect 39564 13582 39566 13634
rect 39618 13582 39620 13634
rect 39564 13524 39620 13582
rect 39564 13458 39620 13468
rect 39900 12962 39956 14364
rect 39900 12910 39902 12962
rect 39954 12910 39956 12962
rect 39900 12898 39956 12910
rect 40012 11732 40068 15148
rect 40460 15092 40628 15148
rect 40124 13746 40180 13758
rect 40124 13694 40126 13746
rect 40178 13694 40180 13746
rect 40124 13636 40180 13694
rect 40124 13570 40180 13580
rect 40348 12964 40404 12974
rect 40348 12870 40404 12908
rect 40012 11676 40180 11732
rect 39452 11508 39508 11518
rect 40012 11508 40068 11518
rect 39452 11506 40068 11508
rect 39452 11454 39454 11506
rect 39506 11454 40014 11506
rect 40066 11454 40068 11506
rect 39452 11452 40068 11454
rect 39452 11442 39508 11452
rect 40012 11442 40068 11452
rect 39340 11228 39508 11284
rect 39340 10724 39396 10734
rect 39228 10722 39396 10724
rect 39228 10670 39342 10722
rect 39394 10670 39396 10722
rect 39228 10668 39396 10670
rect 39340 10658 39396 10668
rect 39116 10558 39118 10610
rect 39170 10558 39172 10610
rect 39116 10546 39172 10558
rect 39452 10612 39508 11228
rect 39900 11282 39956 11294
rect 40124 11284 40180 11676
rect 39900 11230 39902 11282
rect 39954 11230 39956 11282
rect 39900 11060 39956 11230
rect 39900 10994 39956 11004
rect 40012 11228 40180 11284
rect 40236 11396 40292 11406
rect 40460 11396 40516 15092
rect 40572 14644 40628 14654
rect 40572 14530 40628 14588
rect 40572 14478 40574 14530
rect 40626 14478 40628 14530
rect 40572 14466 40628 14478
rect 40684 14306 40740 14318
rect 40684 14254 40686 14306
rect 40738 14254 40740 14306
rect 40684 13524 40740 14254
rect 40908 14308 40964 14318
rect 40908 14306 41188 14308
rect 40908 14254 40910 14306
rect 40962 14254 41188 14306
rect 40908 14252 41188 14254
rect 40908 14242 40964 14252
rect 41020 13524 41076 13534
rect 40684 13468 41020 13524
rect 41020 13430 41076 13468
rect 40236 11394 40516 11396
rect 40236 11342 40238 11394
rect 40290 11342 40516 11394
rect 40236 11340 40516 11342
rect 40012 10722 40068 11228
rect 40236 11172 40292 11340
rect 40236 11106 40292 11116
rect 40684 11172 40740 11182
rect 40684 11078 40740 11116
rect 40012 10670 40014 10722
rect 40066 10670 40068 10722
rect 39564 10612 39620 10622
rect 39452 10610 39620 10612
rect 39452 10558 39566 10610
rect 39618 10558 39620 10610
rect 39452 10556 39620 10558
rect 38780 10388 38836 10398
rect 38780 10386 39284 10388
rect 38780 10334 38782 10386
rect 38834 10334 39284 10386
rect 38780 10332 39284 10334
rect 38780 10322 38836 10332
rect 36428 9874 36484 9884
rect 37660 9996 37828 10052
rect 36428 9714 36484 9726
rect 36428 9662 36430 9714
rect 36482 9662 36484 9714
rect 36428 9604 36484 9662
rect 36428 9538 36484 9548
rect 37100 9604 37156 9614
rect 37100 9154 37156 9548
rect 37100 9102 37102 9154
rect 37154 9102 37156 9154
rect 37100 9090 37156 9102
rect 37212 9154 37268 9166
rect 37212 9102 37214 9154
rect 37266 9102 37268 9154
rect 37212 9044 37268 9102
rect 37212 8988 37604 9044
rect 37212 8820 37268 8830
rect 37212 8818 37380 8820
rect 37212 8766 37214 8818
rect 37266 8766 37380 8818
rect 37212 8764 37380 8766
rect 37212 8754 37268 8764
rect 36979 8652 37243 8662
rect 37035 8596 37083 8652
rect 37139 8596 37187 8652
rect 36979 8586 37243 8596
rect 37212 8484 37268 8494
rect 37324 8484 37380 8764
rect 37212 8482 37380 8484
rect 37212 8430 37214 8482
rect 37266 8430 37380 8482
rect 37212 8428 37380 8430
rect 37548 8484 37604 8988
rect 37212 8418 37268 8428
rect 35868 8206 35870 8258
rect 35922 8206 35924 8258
rect 35868 8194 35924 8206
rect 36092 8372 36148 8382
rect 37436 8372 37492 8382
rect 34076 8082 34132 8092
rect 34972 8148 35028 8158
rect 34972 8054 35028 8092
rect 35532 8148 35588 8158
rect 34524 8036 34580 8046
rect 34188 7588 34244 7598
rect 34076 7532 34188 7588
rect 33964 7252 34020 7262
rect 33964 7158 34020 7196
rect 33740 6692 33796 6702
rect 33292 5966 33294 6018
rect 33346 5966 33348 6018
rect 30828 4338 30996 4340
rect 30828 4286 30830 4338
rect 30882 4286 30996 4338
rect 30828 4284 30996 4286
rect 31164 4340 31220 4350
rect 30828 4274 30884 4284
rect 28924 4162 28980 4172
rect 31164 4226 31220 4284
rect 31164 4174 31166 4226
rect 31218 4174 31220 4226
rect 31164 4162 31220 4174
rect 31948 4338 32004 4350
rect 31948 4286 31950 4338
rect 32002 4286 32004 4338
rect 27356 4114 27524 4116
rect 27356 4062 27358 4114
rect 27410 4062 27524 4114
rect 27356 4060 27524 4062
rect 25676 3668 25732 3678
rect 25676 3574 25732 3612
rect 27356 3668 27412 4060
rect 31948 4004 32004 4286
rect 31948 3938 32004 3948
rect 32172 3668 32228 5068
rect 32396 4452 32452 5852
rect 32508 5684 32564 5694
rect 33068 5684 33124 5694
rect 32508 5682 33124 5684
rect 32508 5630 32510 5682
rect 32562 5630 33070 5682
rect 33122 5630 33124 5682
rect 32508 5628 33124 5630
rect 32508 5618 32564 5628
rect 33068 5618 33124 5628
rect 33292 5460 33348 5966
rect 33628 6578 33684 6590
rect 33628 6526 33630 6578
rect 33682 6526 33684 6578
rect 32844 5404 33348 5460
rect 33404 5684 33460 5694
rect 33628 5684 33684 6526
rect 33740 6578 33796 6636
rect 33964 6692 34020 6702
rect 34076 6692 34132 7532
rect 34188 7494 34244 7532
rect 34524 7474 34580 7980
rect 35084 8036 35140 8046
rect 35084 7942 35140 7980
rect 35420 8036 35476 8046
rect 34860 7700 34916 7710
rect 34860 7698 35252 7700
rect 34860 7646 34862 7698
rect 34914 7646 35252 7698
rect 34860 7644 35252 7646
rect 34860 7634 34916 7644
rect 34524 7422 34526 7474
rect 34578 7422 34580 7474
rect 34524 7410 34580 7422
rect 34748 7476 34804 7486
rect 34748 7382 34804 7420
rect 33964 6690 34132 6692
rect 33964 6638 33966 6690
rect 34018 6638 34132 6690
rect 33964 6636 34132 6638
rect 34636 6692 34692 6702
rect 33964 6626 34020 6636
rect 34636 6598 34692 6636
rect 35196 6692 35252 7644
rect 35420 6802 35476 7980
rect 35532 6916 35588 8092
rect 35644 8034 35700 8046
rect 35644 7982 35646 8034
rect 35698 7982 35700 8034
rect 35644 7588 35700 7982
rect 35644 7522 35700 7532
rect 35644 6916 35700 6926
rect 35532 6914 35700 6916
rect 35532 6862 35646 6914
rect 35698 6862 35700 6914
rect 35532 6860 35700 6862
rect 35420 6750 35422 6802
rect 35474 6750 35476 6802
rect 35420 6692 35476 6750
rect 35196 6690 35364 6692
rect 35196 6638 35198 6690
rect 35250 6638 35364 6690
rect 35196 6636 35364 6638
rect 35196 6626 35252 6636
rect 33740 6526 33742 6578
rect 33794 6526 33796 6578
rect 33740 6514 33796 6526
rect 33404 5682 33684 5684
rect 33404 5630 33406 5682
rect 33458 5630 33684 5682
rect 33404 5628 33684 5630
rect 34972 5906 35028 5918
rect 34972 5854 34974 5906
rect 35026 5854 35028 5906
rect 32508 4452 32564 4462
rect 32396 4450 32564 4452
rect 32396 4398 32510 4450
rect 32562 4398 32564 4450
rect 32396 4396 32564 4398
rect 32508 4386 32564 4396
rect 32284 4340 32340 4350
rect 32284 4246 32340 4284
rect 32284 3668 32340 3678
rect 32172 3666 32676 3668
rect 32172 3614 32286 3666
rect 32338 3614 32676 3666
rect 32172 3612 32676 3614
rect 27356 3602 27412 3612
rect 32284 3602 32340 3612
rect 25564 3556 25620 3566
rect 25508 3554 25620 3556
rect 25508 3502 25566 3554
rect 25618 3502 25620 3554
rect 25508 3500 25620 3502
rect 25452 3462 25508 3500
rect 25564 3490 25620 3500
rect 32620 3554 32676 3612
rect 32844 3666 32900 5404
rect 33404 5236 33460 5628
rect 33404 5170 33460 5180
rect 34412 5236 34468 5246
rect 34412 5142 34468 5180
rect 34524 5236 34580 5246
rect 34860 5236 34916 5246
rect 34972 5236 35028 5854
rect 35196 5908 35252 5918
rect 35196 5814 35252 5852
rect 35084 5796 35140 5806
rect 35084 5702 35140 5740
rect 35084 5348 35140 5358
rect 35308 5348 35364 6636
rect 35420 6626 35476 6636
rect 35644 5906 35700 6860
rect 35644 5854 35646 5906
rect 35698 5854 35700 5906
rect 35644 5842 35700 5854
rect 35756 5908 35812 5918
rect 35084 5346 35364 5348
rect 35084 5294 35086 5346
rect 35138 5294 35364 5346
rect 35084 5292 35364 5294
rect 35756 5346 35812 5852
rect 35756 5294 35758 5346
rect 35810 5294 35812 5346
rect 35084 5282 35140 5292
rect 35756 5282 35812 5294
rect 35868 5684 35924 5694
rect 34524 5234 35028 5236
rect 34524 5182 34526 5234
rect 34578 5182 34862 5234
rect 34914 5182 35028 5234
rect 34524 5180 35028 5182
rect 35868 5234 35924 5628
rect 35868 5182 35870 5234
rect 35922 5182 35924 5234
rect 34524 5170 34580 5180
rect 34860 5170 34916 5180
rect 35868 5170 35924 5182
rect 35420 4898 35476 4910
rect 35420 4846 35422 4898
rect 35474 4846 35476 4898
rect 35420 4788 35476 4846
rect 35420 4722 35476 4732
rect 36092 4788 36148 8316
rect 37324 8370 37492 8372
rect 37324 8318 37438 8370
rect 37490 8318 37492 8370
rect 37324 8316 37492 8318
rect 36979 7084 37243 7094
rect 37035 7028 37083 7084
rect 37139 7028 37187 7084
rect 36979 7018 37243 7028
rect 36092 4722 36148 4732
rect 36316 6692 36372 6702
rect 36316 4562 36372 6636
rect 36988 6132 37044 6142
rect 36988 6038 37044 6076
rect 36979 5516 37243 5526
rect 37035 5460 37083 5516
rect 37139 5460 37187 5516
rect 36979 5450 37243 5460
rect 36876 5012 36932 5022
rect 36316 4510 36318 4562
rect 36370 4510 36372 4562
rect 36316 4498 36372 4510
rect 36764 4956 36876 5012
rect 33292 4450 33348 4462
rect 33292 4398 33294 4450
rect 33346 4398 33348 4450
rect 33068 4340 33124 4350
rect 33068 4246 33124 4284
rect 33180 4226 33236 4238
rect 33180 4174 33182 4226
rect 33234 4174 33236 4226
rect 33180 3892 33236 4174
rect 33292 4004 33348 4398
rect 36652 4116 36708 4126
rect 33292 3938 33348 3948
rect 36540 4114 36708 4116
rect 36540 4062 36654 4114
rect 36706 4062 36708 4114
rect 36540 4060 36708 4062
rect 32956 3836 33236 3892
rect 32956 3778 33012 3836
rect 32956 3726 32958 3778
rect 33010 3726 33012 3778
rect 32956 3714 33012 3726
rect 36540 3778 36596 4060
rect 36652 4050 36708 4060
rect 36540 3726 36542 3778
rect 36594 3726 36596 3778
rect 36540 3714 36596 3726
rect 36764 3780 36820 4956
rect 36876 4946 36932 4956
rect 37324 4450 37380 8316
rect 37436 8306 37492 8316
rect 37436 8148 37492 8158
rect 37548 8148 37604 8428
rect 37436 8146 37604 8148
rect 37436 8094 37438 8146
rect 37490 8094 37604 8146
rect 37436 8092 37604 8094
rect 37436 8082 37492 8092
rect 37548 6132 37604 6142
rect 37660 6132 37716 9996
rect 38444 9940 38500 9950
rect 38444 9846 38500 9884
rect 37772 9828 37828 9838
rect 37772 8370 37828 9772
rect 38108 9826 38164 9838
rect 38108 9774 38110 9826
rect 38162 9774 38164 9826
rect 38108 9716 38164 9774
rect 38332 9716 38388 9726
rect 38164 9660 38276 9716
rect 38108 9650 38164 9660
rect 37772 8318 37774 8370
rect 37826 8318 37828 8370
rect 37772 8306 37828 8318
rect 37996 8260 38052 8270
rect 38108 8260 38164 8270
rect 37996 8258 38108 8260
rect 37996 8206 37998 8258
rect 38050 8206 38108 8258
rect 37996 8204 38108 8206
rect 37996 8194 38052 8204
rect 37604 6076 37716 6132
rect 37548 6038 37604 6076
rect 37660 5460 37716 6076
rect 37884 5908 37940 5918
rect 37884 5814 37940 5852
rect 37660 5234 37716 5404
rect 37660 5182 37662 5234
rect 37714 5182 37716 5234
rect 37660 5170 37716 5182
rect 37996 4898 38052 4910
rect 37996 4846 37998 4898
rect 38050 4846 38052 4898
rect 37324 4398 37326 4450
rect 37378 4398 37380 4450
rect 37324 4386 37380 4398
rect 37436 4676 37492 4686
rect 37436 4338 37492 4620
rect 37436 4286 37438 4338
rect 37490 4286 37492 4338
rect 37436 4274 37492 4286
rect 36979 3948 37243 3958
rect 37035 3892 37083 3948
rect 37139 3892 37187 3948
rect 36979 3882 37243 3892
rect 36876 3780 36932 3790
rect 36764 3778 36932 3780
rect 36764 3726 36878 3778
rect 36930 3726 36932 3778
rect 36764 3724 36932 3726
rect 36876 3714 36932 3724
rect 32844 3614 32846 3666
rect 32898 3614 32900 3666
rect 32844 3602 32900 3614
rect 32620 3502 32622 3554
rect 32674 3502 32676 3554
rect 32620 3490 32676 3502
rect 37548 3556 37604 3566
rect 24668 3390 24670 3442
rect 24722 3390 24724 3442
rect 24668 3378 24724 3390
rect 25788 3444 25844 3482
rect 37548 3462 37604 3500
rect 25788 3378 25844 3388
rect 37660 3444 37716 3454
rect 37996 3444 38052 4846
rect 38108 3556 38164 8204
rect 38220 6916 38276 9660
rect 38332 9622 38388 9660
rect 39228 8708 39284 10332
rect 39340 9716 39396 9726
rect 39340 9622 39396 9660
rect 39452 9268 39508 9278
rect 39452 9174 39508 9212
rect 39228 8652 39396 8708
rect 39228 8482 39284 8494
rect 39228 8430 39230 8482
rect 39282 8430 39284 8482
rect 39228 8260 39284 8430
rect 39228 8194 39284 8204
rect 39340 8258 39396 8652
rect 39340 8206 39342 8258
rect 39394 8206 39396 8258
rect 39340 8036 39396 8206
rect 38780 7980 39396 8036
rect 38780 7586 38836 7980
rect 38780 7534 38782 7586
rect 38834 7534 38836 7586
rect 38220 6860 38388 6916
rect 38220 6690 38276 6702
rect 38220 6638 38222 6690
rect 38274 6638 38276 6690
rect 38220 6130 38276 6638
rect 38220 6078 38222 6130
rect 38274 6078 38276 6130
rect 38220 6066 38276 6078
rect 38332 5908 38388 6860
rect 38780 6580 38836 7534
rect 39116 7250 39172 7262
rect 39116 7198 39118 7250
rect 39170 7198 39172 7250
rect 38220 5906 38388 5908
rect 38220 5854 38334 5906
rect 38386 5854 38388 5906
rect 38220 5852 38388 5854
rect 38220 5012 38276 5852
rect 38332 5842 38388 5852
rect 38444 6524 38836 6580
rect 39004 6580 39060 6590
rect 38444 6018 38500 6524
rect 39004 6486 39060 6524
rect 39116 6356 39172 7198
rect 39228 6692 39284 6702
rect 39564 6692 39620 10556
rect 39788 10498 39844 10510
rect 39788 10446 39790 10498
rect 39842 10446 39844 10498
rect 39788 9940 39844 10446
rect 39788 9874 39844 9884
rect 40012 9268 40068 10670
rect 40124 10836 40180 10846
rect 40124 10610 40180 10780
rect 41132 10724 41188 14252
rect 41244 13972 41300 15260
rect 41244 13906 41300 13916
rect 41356 14530 41412 15484
rect 41468 14642 41524 16492
rect 41692 16210 41748 16716
rect 41692 16158 41694 16210
rect 41746 16158 41748 16210
rect 41692 16146 41748 16158
rect 42140 15540 42196 15550
rect 42140 15446 42196 15484
rect 42588 15538 42644 16828
rect 43484 16882 43540 17052
rect 43596 16994 43652 17164
rect 43932 17108 43988 18396
rect 44132 17276 44396 17286
rect 44188 17220 44236 17276
rect 44292 17220 44340 17276
rect 44132 17210 44396 17220
rect 43932 17052 44324 17108
rect 43596 16942 43598 16994
rect 43650 16942 43652 16994
rect 43596 16930 43652 16942
rect 44268 16994 44324 17052
rect 44268 16942 44270 16994
rect 44322 16942 44324 16994
rect 44268 16930 44324 16942
rect 43484 16830 43486 16882
rect 43538 16830 43540 16882
rect 43484 16818 43540 16830
rect 43708 16772 43764 16782
rect 44156 16772 44212 16782
rect 43708 16098 43764 16716
rect 43708 16046 43710 16098
rect 43762 16046 43764 16098
rect 43708 16034 43764 16046
rect 43932 16770 44212 16772
rect 43932 16718 44158 16770
rect 44210 16718 44212 16770
rect 43932 16716 44212 16718
rect 43932 16100 43988 16716
rect 44156 16706 44212 16716
rect 44492 16436 44548 18956
rect 44716 18564 44772 18574
rect 44828 18564 44884 22316
rect 45948 22370 46004 22382
rect 45948 22318 45950 22370
rect 46002 22318 46004 22370
rect 45276 22260 45332 22270
rect 45276 21698 45332 22204
rect 45948 21700 46004 22318
rect 45276 21646 45278 21698
rect 45330 21646 45332 21698
rect 45276 21634 45332 21646
rect 45836 21644 45948 21700
rect 45052 21362 45108 21374
rect 45052 21310 45054 21362
rect 45106 21310 45108 21362
rect 44940 20580 44996 20590
rect 44940 19908 44996 20524
rect 45052 20130 45108 21310
rect 45836 20802 45892 21644
rect 45948 21634 46004 21644
rect 46060 22258 46116 22270
rect 46060 22206 46062 22258
rect 46114 22206 46116 22258
rect 45836 20750 45838 20802
rect 45890 20750 45892 20802
rect 45836 20244 45892 20750
rect 46060 20804 46116 22206
rect 46060 20710 46116 20748
rect 45836 20178 45892 20188
rect 45052 20078 45054 20130
rect 45106 20078 45108 20130
rect 45052 20066 45108 20078
rect 45948 20132 46004 20142
rect 44940 19852 45108 19908
rect 45052 19458 45108 19852
rect 45276 19796 45332 19806
rect 45052 19406 45054 19458
rect 45106 19406 45108 19458
rect 45052 19394 45108 19406
rect 45164 19740 45276 19796
rect 45164 19236 45220 19740
rect 45276 19730 45332 19740
rect 45948 19460 46004 20076
rect 46284 20020 46340 23662
rect 46508 23154 46564 23166
rect 46508 23102 46510 23154
rect 46562 23102 46564 23154
rect 46508 22484 46564 23102
rect 47068 23156 47124 23774
rect 47180 23828 47236 23886
rect 47180 23762 47236 23772
rect 47068 23062 47124 23100
rect 47292 23266 47348 23278
rect 47292 23214 47294 23266
rect 47346 23214 47348 23266
rect 46956 23042 47012 23054
rect 46956 22990 46958 23042
rect 47010 22990 47012 23042
rect 46956 22596 47012 22990
rect 46508 21924 46564 22428
rect 46508 21858 46564 21868
rect 46844 22540 46956 22596
rect 46284 19926 46340 19964
rect 46620 21586 46676 21598
rect 46620 21534 46622 21586
rect 46674 21534 46676 21586
rect 46620 21476 46676 21534
rect 46172 19796 46228 19806
rect 46172 19702 46228 19740
rect 45500 19458 46004 19460
rect 45500 19406 45950 19458
rect 46002 19406 46004 19458
rect 45500 19404 46004 19406
rect 44716 18562 44884 18564
rect 44716 18510 44718 18562
rect 44770 18510 44884 18562
rect 44716 18508 44884 18510
rect 45052 19180 45220 19236
rect 45276 19236 45332 19246
rect 44604 18340 44660 18350
rect 44604 16882 44660 18284
rect 44716 17668 44772 18508
rect 44716 17602 44772 17612
rect 45052 17666 45108 19180
rect 45276 19122 45332 19180
rect 45276 19070 45278 19122
rect 45330 19070 45332 19122
rect 45276 19058 45332 19070
rect 45164 19012 45220 19022
rect 45164 18918 45220 18956
rect 45052 17614 45054 17666
rect 45106 17614 45108 17666
rect 45052 17602 45108 17614
rect 45164 18674 45220 18686
rect 45164 18622 45166 18674
rect 45218 18622 45220 18674
rect 44604 16830 44606 16882
rect 44658 16830 44660 16882
rect 44604 16818 44660 16830
rect 43932 16006 43988 16044
rect 44268 16380 44548 16436
rect 43820 15876 43876 15886
rect 44268 15876 44324 16380
rect 45164 16324 45220 18622
rect 45500 18450 45556 19404
rect 45948 19394 46004 19404
rect 46060 19684 46116 19694
rect 46060 19234 46116 19628
rect 46060 19182 46062 19234
rect 46114 19182 46116 19234
rect 46060 19170 46116 19182
rect 46508 19572 46564 19582
rect 46396 18452 46452 18462
rect 45500 18398 45502 18450
rect 45554 18398 45556 18450
rect 45500 18386 45556 18398
rect 45612 18450 46452 18452
rect 45612 18398 46398 18450
rect 46450 18398 46452 18450
rect 45612 18396 46452 18398
rect 45276 18116 45332 18126
rect 45276 17778 45332 18060
rect 45276 17726 45278 17778
rect 45330 17726 45332 17778
rect 45276 17714 45332 17726
rect 45612 17778 45668 18396
rect 46396 18386 46452 18396
rect 46508 18228 46564 19516
rect 46620 19236 46676 21420
rect 46732 20804 46788 20814
rect 46732 19460 46788 20748
rect 46844 19684 46900 22540
rect 46956 22530 47012 22540
rect 47068 22372 47124 22382
rect 47068 22278 47124 22316
rect 47292 22372 47348 23214
rect 46956 22148 47012 22158
rect 47292 22148 47348 22316
rect 46956 22146 47348 22148
rect 46956 22094 46958 22146
rect 47010 22094 47348 22146
rect 46956 22092 47348 22094
rect 46956 22082 47012 22092
rect 47628 22036 47684 24668
rect 48188 24612 48244 24622
rect 48188 24518 48244 24556
rect 48076 24498 48132 24510
rect 48076 24446 48078 24498
rect 48130 24446 48132 24498
rect 47964 22260 48020 22270
rect 47964 22166 48020 22204
rect 47516 21980 47684 22036
rect 47740 22148 47796 22158
rect 47404 21698 47460 21710
rect 47404 21646 47406 21698
rect 47458 21646 47460 21698
rect 47180 21586 47236 21598
rect 47180 21534 47182 21586
rect 47234 21534 47236 21586
rect 47180 21028 47236 21534
rect 47404 21476 47460 21646
rect 47180 20962 47236 20972
rect 47292 21420 47404 21476
rect 46844 19618 46900 19628
rect 46956 20690 47012 20702
rect 46956 20638 46958 20690
rect 47010 20638 47012 20690
rect 46956 20020 47012 20638
rect 47068 20132 47124 20142
rect 47068 20038 47124 20076
rect 46732 19394 46788 19404
rect 46956 19236 47012 19964
rect 46620 19180 46900 19236
rect 46732 18452 46788 18462
rect 46732 18358 46788 18396
rect 46844 18452 46900 19180
rect 46956 19170 47012 19180
rect 47180 19908 47236 19918
rect 47068 18452 47124 18462
rect 46844 18450 47124 18452
rect 46844 18398 47070 18450
rect 47122 18398 47124 18450
rect 46844 18396 47124 18398
rect 46844 18340 46900 18396
rect 47068 18386 47124 18396
rect 46844 18274 46900 18284
rect 45612 17726 45614 17778
rect 45666 17726 45668 17778
rect 45612 17714 45668 17726
rect 46396 18172 46564 18228
rect 46284 17668 46340 17678
rect 46284 17574 46340 17612
rect 45388 17108 45444 17118
rect 45388 17014 45444 17052
rect 44380 16268 45220 16324
rect 44380 16098 44436 16268
rect 45164 16210 45220 16268
rect 45164 16158 45166 16210
rect 45218 16158 45220 16210
rect 45164 16146 45220 16158
rect 44380 16046 44382 16098
rect 44434 16046 44436 16098
rect 44380 16034 44436 16046
rect 45052 16100 45108 16110
rect 45052 16006 45108 16044
rect 45836 15988 45892 15998
rect 45724 15876 45780 15886
rect 44268 15820 44884 15876
rect 43820 15782 43876 15820
rect 44132 15708 44396 15718
rect 44188 15652 44236 15708
rect 44292 15652 44340 15708
rect 44132 15642 44396 15652
rect 42588 15486 42590 15538
rect 42642 15486 42644 15538
rect 42588 15474 42644 15486
rect 44604 15540 44660 15550
rect 44604 15446 44660 15484
rect 44828 15538 44884 15820
rect 44828 15486 44830 15538
rect 44882 15486 44884 15538
rect 41692 15426 41748 15438
rect 41692 15374 41694 15426
rect 41746 15374 41748 15426
rect 41580 15316 41636 15326
rect 41580 15202 41636 15260
rect 41580 15150 41582 15202
rect 41634 15150 41636 15202
rect 41580 15138 41636 15150
rect 41468 14590 41470 14642
rect 41522 14590 41524 14642
rect 41468 14578 41524 14590
rect 41692 14532 41748 15374
rect 42364 15316 42420 15326
rect 42364 15222 42420 15260
rect 44268 15314 44324 15326
rect 44268 15262 44270 15314
rect 44322 15262 44324 15314
rect 41356 14478 41358 14530
rect 41410 14478 41412 14530
rect 41356 13746 41412 14478
rect 41580 14530 41748 14532
rect 41580 14478 41694 14530
rect 41746 14478 41748 14530
rect 41580 14476 41748 14478
rect 41580 13860 41636 14476
rect 41692 14466 41748 14476
rect 42476 15202 42532 15214
rect 42476 15150 42478 15202
rect 42530 15150 42532 15202
rect 41916 14306 41972 14318
rect 41916 14254 41918 14306
rect 41970 14254 41972 14306
rect 41580 13766 41636 13804
rect 41692 13972 41748 13982
rect 41356 13694 41358 13746
rect 41410 13694 41412 13746
rect 41356 13682 41412 13694
rect 41244 13636 41300 13646
rect 41244 12850 41300 13580
rect 41244 12798 41246 12850
rect 41298 12798 41300 12850
rect 41244 12786 41300 12798
rect 41356 12738 41412 12750
rect 41356 12686 41358 12738
rect 41410 12686 41412 12738
rect 41244 10724 41300 10734
rect 41132 10722 41300 10724
rect 41132 10670 41246 10722
rect 41298 10670 41300 10722
rect 41132 10668 41300 10670
rect 40124 10558 40126 10610
rect 40178 10558 40180 10610
rect 40124 10546 40180 10558
rect 40908 10498 40964 10510
rect 40908 10446 40910 10498
rect 40962 10446 40964 10498
rect 40348 10164 40404 10174
rect 40124 9940 40180 9950
rect 40348 9940 40404 10108
rect 40348 9884 40516 9940
rect 40124 9826 40180 9884
rect 40124 9774 40126 9826
rect 40178 9774 40180 9826
rect 40124 9762 40180 9774
rect 40460 9826 40516 9884
rect 40460 9774 40462 9826
rect 40514 9774 40516 9826
rect 40348 9716 40404 9726
rect 40012 9202 40068 9212
rect 40236 9714 40404 9716
rect 40236 9662 40350 9714
rect 40402 9662 40404 9714
rect 40236 9660 40404 9662
rect 40236 8932 40292 9660
rect 40348 9650 40404 9660
rect 40460 9156 40516 9774
rect 40908 9716 40964 10446
rect 41244 10052 41300 10668
rect 41244 9986 41300 9996
rect 40908 9380 40964 9660
rect 40460 9090 40516 9100
rect 40572 9324 40964 9380
rect 40124 7476 40180 7486
rect 40124 7382 40180 7420
rect 39228 6690 39620 6692
rect 39228 6638 39230 6690
rect 39282 6638 39620 6690
rect 39228 6636 39620 6638
rect 40124 6692 40180 6702
rect 39228 6626 39284 6636
rect 39004 6300 39172 6356
rect 38444 5966 38446 6018
rect 38498 5966 38500 6018
rect 38332 5460 38388 5470
rect 38332 5346 38388 5404
rect 38332 5294 38334 5346
rect 38386 5294 38388 5346
rect 38332 5282 38388 5294
rect 38444 5236 38500 5966
rect 38444 5170 38500 5180
rect 38556 6244 38612 6254
rect 38556 5234 38612 6188
rect 38556 5182 38558 5234
rect 38610 5182 38612 5234
rect 38556 5170 38612 5182
rect 39004 6244 39060 6300
rect 38220 4946 38276 4956
rect 38668 5124 38724 5134
rect 38668 4450 38724 5068
rect 38668 4398 38670 4450
rect 38722 4398 38724 4450
rect 38668 4386 38724 4398
rect 39004 4226 39060 6188
rect 39900 6132 39956 6142
rect 39452 5908 39508 5918
rect 39788 5908 39844 5918
rect 39508 5906 39844 5908
rect 39508 5854 39790 5906
rect 39842 5854 39844 5906
rect 39508 5852 39844 5854
rect 39228 5236 39284 5246
rect 39116 4900 39172 4910
rect 39116 4806 39172 4844
rect 39228 4900 39284 5180
rect 39452 5124 39508 5852
rect 39788 5842 39844 5852
rect 39900 5684 39956 6076
rect 40124 6130 40180 6636
rect 40236 6244 40292 8876
rect 40572 8484 40628 9324
rect 41020 9268 41076 9278
rect 40572 8418 40628 8428
rect 40684 9266 41076 9268
rect 40684 9214 41022 9266
rect 41074 9214 41076 9266
rect 40684 9212 41076 9214
rect 40684 8258 40740 9212
rect 41020 9202 41076 9212
rect 40908 9044 40964 9054
rect 40684 8206 40686 8258
rect 40738 8206 40740 8258
rect 40684 8194 40740 8206
rect 40796 8484 40852 8494
rect 40796 6692 40852 8428
rect 40908 7586 40964 8988
rect 41132 9044 41188 9054
rect 41356 9044 41412 12686
rect 41692 11620 41748 13916
rect 41580 11564 41748 11620
rect 41804 12178 41860 12190
rect 41804 12126 41806 12178
rect 41858 12126 41860 12178
rect 41580 10612 41636 11564
rect 41692 11396 41748 11406
rect 41804 11396 41860 12126
rect 41916 12068 41972 14254
rect 42028 13748 42084 13758
rect 42028 13654 42084 13692
rect 42252 13746 42308 13758
rect 42252 13694 42254 13746
rect 42306 13694 42308 13746
rect 42252 13524 42308 13694
rect 42252 13458 42308 13468
rect 42028 12068 42084 12078
rect 41916 12066 42084 12068
rect 41916 12014 42030 12066
rect 42082 12014 42084 12066
rect 41916 12012 42084 12014
rect 41916 11506 41972 12012
rect 42028 12002 42084 12012
rect 41916 11454 41918 11506
rect 41970 11454 41972 11506
rect 41916 11442 41972 11454
rect 41692 11394 41860 11396
rect 41692 11342 41694 11394
rect 41746 11342 41860 11394
rect 41692 11340 41860 11342
rect 41692 11060 41748 11340
rect 41692 10994 41748 11004
rect 42028 10722 42084 10734
rect 42028 10670 42030 10722
rect 42082 10670 42084 10722
rect 41916 10612 41972 10622
rect 41580 10610 41748 10612
rect 41580 10558 41582 10610
rect 41634 10558 41748 10610
rect 41580 10556 41748 10558
rect 41580 10546 41636 10556
rect 41580 9156 41636 9166
rect 41580 9062 41636 9100
rect 41132 9042 41412 9044
rect 41132 8990 41134 9042
rect 41186 8990 41412 9042
rect 41132 8988 41412 8990
rect 41020 8372 41076 8382
rect 41020 7698 41076 8316
rect 41020 7646 41022 7698
rect 41074 7646 41076 7698
rect 41020 7634 41076 7646
rect 40908 7534 40910 7586
rect 40962 7534 40964 7586
rect 40908 7522 40964 7534
rect 41132 7476 41188 8988
rect 41692 8372 41748 10556
rect 41692 8306 41748 8316
rect 41804 9938 41860 9950
rect 41804 9886 41806 9938
rect 41858 9886 41860 9938
rect 41804 8260 41860 9886
rect 41916 9042 41972 10556
rect 42028 9156 42084 10670
rect 42252 10610 42308 10622
rect 42252 10558 42254 10610
rect 42306 10558 42308 10610
rect 42028 9090 42084 9100
rect 42140 10052 42196 10062
rect 41916 8990 41918 9042
rect 41970 8990 41972 9042
rect 41916 8484 41972 8990
rect 41916 8428 42084 8484
rect 41804 8166 41860 8204
rect 42028 8148 42084 8428
rect 42140 8370 42196 9996
rect 42252 9380 42308 10558
rect 42476 9828 42532 15150
rect 42700 14756 42756 14766
rect 42700 12404 42756 14700
rect 44268 14532 44324 15262
rect 44828 15148 44884 15486
rect 45388 15540 45444 15550
rect 45388 15446 45444 15484
rect 45724 15426 45780 15820
rect 45836 15538 45892 15932
rect 45836 15486 45838 15538
rect 45890 15486 45892 15538
rect 45836 15474 45892 15486
rect 45724 15374 45726 15426
rect 45778 15374 45780 15426
rect 45724 15362 45780 15374
rect 46396 15148 46452 18172
rect 47180 16994 47236 19852
rect 47292 19234 47348 21420
rect 47404 21410 47460 21420
rect 47404 20802 47460 20814
rect 47404 20750 47406 20802
rect 47458 20750 47460 20802
rect 47404 20580 47460 20750
rect 47404 20514 47460 20524
rect 47516 20356 47572 21980
rect 47628 21812 47684 21822
rect 47628 21474 47684 21756
rect 47628 21422 47630 21474
rect 47682 21422 47684 21474
rect 47628 21410 47684 21422
rect 47404 20300 47572 20356
rect 47404 19572 47460 20300
rect 47404 19506 47460 19516
rect 47516 20132 47572 20142
rect 47292 19182 47294 19234
rect 47346 19182 47348 19234
rect 47292 19170 47348 19182
rect 47180 16942 47182 16994
rect 47234 16942 47236 16994
rect 47180 16930 47236 16942
rect 47516 16994 47572 20076
rect 47740 20018 47796 22092
rect 48076 20916 48132 24446
rect 48636 23940 48692 23950
rect 48972 23940 49028 25228
rect 49084 24722 49140 26798
rect 49756 26850 49812 26862
rect 49756 26798 49758 26850
rect 49810 26798 49812 26850
rect 49756 26402 49812 26798
rect 50316 26516 50372 27244
rect 50316 26422 50372 26460
rect 52220 26516 52276 26526
rect 52220 26422 52276 26460
rect 57708 26514 57764 27356
rect 58439 26684 58703 26694
rect 58495 26628 58543 26684
rect 58599 26628 58647 26684
rect 58439 26618 58703 26628
rect 57708 26462 57710 26514
rect 57762 26462 57764 26514
rect 57708 26450 57764 26462
rect 49756 26350 49758 26402
rect 49810 26350 49812 26402
rect 49756 26338 49812 26350
rect 50652 26402 50708 26414
rect 50652 26350 50654 26402
rect 50706 26350 50708 26402
rect 49532 26292 49588 26302
rect 49196 26068 49252 26078
rect 49196 25974 49252 26012
rect 49196 25396 49252 25406
rect 49532 25396 49588 26236
rect 49980 26292 50036 26302
rect 49980 26198 50036 26236
rect 50428 26292 50484 26302
rect 50204 26068 50260 26078
rect 50428 26068 50484 26236
rect 50260 26012 50372 26068
rect 50204 26002 50260 26012
rect 49252 25340 49700 25396
rect 49196 25302 49252 25340
rect 49084 24670 49086 24722
rect 49138 24670 49140 24722
rect 49084 24658 49140 24670
rect 49196 24946 49252 24958
rect 49196 24894 49198 24946
rect 49250 24894 49252 24946
rect 49196 24612 49252 24894
rect 49644 24834 49700 25340
rect 49644 24782 49646 24834
rect 49698 24782 49700 24834
rect 49644 24770 49700 24782
rect 50204 25282 50260 25294
rect 50204 25230 50206 25282
rect 50258 25230 50260 25282
rect 49196 24556 50036 24612
rect 49532 23940 49588 23950
rect 48972 23938 49588 23940
rect 48972 23886 49534 23938
rect 49586 23886 49588 23938
rect 48972 23884 49588 23886
rect 48636 23826 48692 23884
rect 48636 23774 48638 23826
rect 48690 23774 48692 23826
rect 48636 23762 48692 23774
rect 48748 23828 48804 23838
rect 48412 23156 48468 23166
rect 48412 22370 48468 23100
rect 48412 22318 48414 22370
rect 48466 22318 48468 22370
rect 48412 22306 48468 22318
rect 48748 23154 48804 23772
rect 49532 23268 49588 23884
rect 49532 23174 49588 23212
rect 49644 23826 49700 23838
rect 49644 23774 49646 23826
rect 49698 23774 49700 23826
rect 48748 23102 48750 23154
rect 48802 23102 48804 23154
rect 48748 22484 48804 23102
rect 48748 21812 48804 22428
rect 49420 22594 49476 22606
rect 49420 22542 49422 22594
rect 49474 22542 49476 22594
rect 48524 21756 48804 21812
rect 48972 22036 49028 22046
rect 48188 21476 48244 21486
rect 48188 21382 48244 21420
rect 48076 20914 48244 20916
rect 48076 20862 48078 20914
rect 48130 20862 48244 20914
rect 48076 20860 48244 20862
rect 48076 20850 48132 20860
rect 47964 20580 48020 20590
rect 47740 19966 47742 20018
rect 47794 19966 47796 20018
rect 47740 19954 47796 19966
rect 47852 20524 47964 20580
rect 47628 18452 47684 18462
rect 47628 17666 47684 18396
rect 47628 17614 47630 17666
rect 47682 17614 47684 17666
rect 47628 17602 47684 17614
rect 47516 16942 47518 16994
rect 47570 16942 47572 16994
rect 47516 16930 47572 16942
rect 47740 16772 47796 16782
rect 47852 16772 47908 20524
rect 47964 20514 48020 20524
rect 48076 20468 48132 20478
rect 48076 20020 48132 20412
rect 47964 19964 48132 20020
rect 47964 19234 48020 19964
rect 47964 19182 47966 19234
rect 48018 19182 48020 19234
rect 47964 19170 48020 19182
rect 48076 19794 48132 19806
rect 48076 19742 48078 19794
rect 48130 19742 48132 19794
rect 48076 18452 48132 19742
rect 48188 18564 48244 20860
rect 48524 20802 48580 21756
rect 48748 21588 48804 21598
rect 48748 21494 48804 21532
rect 48972 21586 49028 21980
rect 49308 21700 49364 21710
rect 49308 21606 49364 21644
rect 48972 21534 48974 21586
rect 49026 21534 49028 21586
rect 48972 21522 49028 21534
rect 48524 20750 48526 20802
rect 48578 20750 48580 20802
rect 48524 20738 48580 20750
rect 48636 21476 48692 21486
rect 48636 20132 48692 21420
rect 48860 20692 48916 20702
rect 49196 20692 49252 20702
rect 48860 20690 49252 20692
rect 48860 20638 48862 20690
rect 48914 20638 49198 20690
rect 49250 20638 49252 20690
rect 48860 20636 49252 20638
rect 48860 20626 48916 20636
rect 49196 20626 49252 20636
rect 49420 20244 49476 22542
rect 49532 22372 49588 22382
rect 49532 22278 49588 22316
rect 49532 21924 49588 21934
rect 49532 20802 49588 21868
rect 49532 20750 49534 20802
rect 49586 20750 49588 20802
rect 49532 20738 49588 20750
rect 49644 21812 49700 23774
rect 49420 20188 49588 20244
rect 49196 20132 49252 20142
rect 48636 20130 49252 20132
rect 48636 20078 49198 20130
rect 49250 20078 49252 20130
rect 48636 20076 49252 20078
rect 48972 19906 49028 19918
rect 48972 19854 48974 19906
rect 49026 19854 49028 19906
rect 48188 18498 48244 18508
rect 48748 19794 48804 19806
rect 48748 19742 48750 19794
rect 48802 19742 48804 19794
rect 48076 18386 48132 18396
rect 48748 18228 48804 19742
rect 48972 19684 49028 19854
rect 48972 19618 49028 19628
rect 49196 19460 49252 20076
rect 49420 20020 49476 20030
rect 49308 19908 49364 19918
rect 49308 19814 49364 19852
rect 49196 19404 49364 19460
rect 49196 19234 49252 19246
rect 49196 19182 49198 19234
rect 49250 19182 49252 19234
rect 49196 19122 49252 19182
rect 49196 19070 49198 19122
rect 49250 19070 49252 19122
rect 49196 19058 49252 19070
rect 48860 18564 48916 18574
rect 48860 18470 48916 18508
rect 49196 18450 49252 18462
rect 49196 18398 49198 18450
rect 49250 18398 49252 18450
rect 49196 18340 49252 18398
rect 49196 18274 49252 18284
rect 48300 17668 48356 17678
rect 48076 17666 48356 17668
rect 48076 17614 48302 17666
rect 48354 17614 48356 17666
rect 48076 17612 48356 17614
rect 48076 17106 48132 17612
rect 48300 17602 48356 17612
rect 48076 17054 48078 17106
rect 48130 17054 48132 17106
rect 48076 17042 48132 17054
rect 48748 17108 48804 18172
rect 48860 17108 48916 17118
rect 48748 17106 48916 17108
rect 48748 17054 48862 17106
rect 48914 17054 48916 17106
rect 48748 17052 48916 17054
rect 48860 17042 48916 17052
rect 49308 17108 49364 19404
rect 49420 19122 49476 19964
rect 49420 19070 49422 19122
rect 49474 19070 49476 19122
rect 49420 19058 49476 19070
rect 49420 18564 49476 18574
rect 49420 17554 49476 18508
rect 49532 18340 49588 20188
rect 49644 19346 49700 21756
rect 49644 19294 49646 19346
rect 49698 19294 49700 19346
rect 49644 19282 49700 19294
rect 49756 23268 49812 23278
rect 49756 22260 49812 23212
rect 49756 19010 49812 22204
rect 49868 19236 49924 19246
rect 49868 19142 49924 19180
rect 49756 18958 49758 19010
rect 49810 18958 49812 19010
rect 49756 18946 49812 18958
rect 49532 18274 49588 18284
rect 49756 18676 49812 18686
rect 49420 17502 49422 17554
rect 49474 17502 49476 17554
rect 49420 17490 49476 17502
rect 49756 17554 49812 18620
rect 49756 17502 49758 17554
rect 49810 17502 49812 17554
rect 49756 17490 49812 17502
rect 49308 17014 49364 17052
rect 47740 16770 47908 16772
rect 47740 16718 47742 16770
rect 47794 16718 47908 16770
rect 47740 16716 47908 16718
rect 47740 16706 47796 16716
rect 47628 16098 47684 16110
rect 47628 16046 47630 16098
rect 47682 16046 47684 16098
rect 46508 15988 46564 15998
rect 46508 15894 46564 15932
rect 47628 15988 47684 16046
rect 47628 15922 47684 15932
rect 47852 16098 47908 16110
rect 47852 16046 47854 16098
rect 47906 16046 47908 16098
rect 47852 15428 47908 16046
rect 48972 16100 49028 16110
rect 47964 15988 48020 15998
rect 47964 15540 48020 15932
rect 48076 15988 48132 15998
rect 48076 15986 48468 15988
rect 48076 15934 48078 15986
rect 48130 15934 48468 15986
rect 48076 15932 48468 15934
rect 48076 15922 48132 15932
rect 48076 15540 48132 15550
rect 47964 15538 48132 15540
rect 47964 15486 48078 15538
rect 48130 15486 48132 15538
rect 47964 15484 48132 15486
rect 48076 15474 48132 15484
rect 47852 15334 47908 15372
rect 47516 15316 47572 15326
rect 44268 14466 44324 14476
rect 44492 15090 44548 15102
rect 44828 15092 45108 15148
rect 44492 15038 44494 15090
rect 44546 15038 44548 15090
rect 44492 14420 44548 15038
rect 44828 14532 44884 14542
rect 44828 14438 44884 14476
rect 45052 14530 45108 15092
rect 45052 14478 45054 14530
rect 45106 14478 45108 14530
rect 45052 14466 45108 14478
rect 45836 15090 45892 15102
rect 45836 15038 45838 15090
rect 45890 15038 45892 15090
rect 44604 14420 44660 14430
rect 44492 14364 44604 14420
rect 44604 14354 44660 14364
rect 45276 14420 45332 14430
rect 45276 14326 45332 14364
rect 45836 14420 45892 15038
rect 45836 14354 45892 14364
rect 46172 15092 46452 15148
rect 47404 15260 47516 15316
rect 44940 14306 44996 14318
rect 44940 14254 44942 14306
rect 44994 14254 44996 14306
rect 44132 14140 44396 14150
rect 44188 14084 44236 14140
rect 44292 14084 44340 14140
rect 44132 14074 44396 14084
rect 44940 13972 44996 14254
rect 45052 13972 45108 13982
rect 44940 13970 45108 13972
rect 44940 13918 45054 13970
rect 45106 13918 45108 13970
rect 44940 13916 45108 13918
rect 45052 13906 45108 13916
rect 44604 13860 44660 13870
rect 44604 13766 44660 13804
rect 45500 13860 45556 13870
rect 45500 13766 45556 13804
rect 44828 13746 44884 13758
rect 44828 13694 44830 13746
rect 44882 13694 44884 13746
rect 42700 12338 42756 12348
rect 42924 13634 42980 13646
rect 42924 13582 42926 13634
rect 42978 13582 42980 13634
rect 42924 11844 42980 13582
rect 44156 13636 44212 13646
rect 44828 13636 44884 13694
rect 45724 13748 45780 13758
rect 45724 13654 45780 13692
rect 44156 13634 44884 13636
rect 44156 13582 44158 13634
rect 44210 13582 44884 13634
rect 44156 13580 44884 13582
rect 44940 13634 44996 13646
rect 44940 13582 44942 13634
rect 44994 13582 44996 13634
rect 44156 12740 44212 13580
rect 44940 12964 44996 13582
rect 45388 13522 45444 13534
rect 45388 13470 45390 13522
rect 45442 13470 45444 13522
rect 45388 13300 45444 13470
rect 45164 13244 45444 13300
rect 45164 13076 45220 13244
rect 46172 13186 46228 15092
rect 46172 13134 46174 13186
rect 46226 13134 46228 13186
rect 46172 13122 46228 13134
rect 46732 13188 46788 13198
rect 45164 12982 45220 13020
rect 46732 13074 46788 13132
rect 46732 13022 46734 13074
rect 46786 13022 46788 13074
rect 46732 13010 46788 13022
rect 47292 13188 47348 13198
rect 44940 12898 44996 12908
rect 45500 12964 45556 12974
rect 45500 12870 45556 12908
rect 43932 12684 44212 12740
rect 45836 12740 45892 12750
rect 46060 12740 46116 12750
rect 42924 11778 42980 11788
rect 43036 12066 43092 12078
rect 43036 12014 43038 12066
rect 43090 12014 43092 12066
rect 42924 11170 42980 11182
rect 42924 11118 42926 11170
rect 42978 11118 42980 11170
rect 42924 10164 42980 11118
rect 43036 10612 43092 12014
rect 43932 11284 43988 12684
rect 45836 12646 45892 12684
rect 45948 12738 46116 12740
rect 45948 12686 46062 12738
rect 46114 12686 46116 12738
rect 45948 12684 46116 12686
rect 44132 12572 44396 12582
rect 44188 12516 44236 12572
rect 44292 12516 44340 12572
rect 45948 12516 46004 12684
rect 46060 12674 46116 12684
rect 47068 12740 47124 12750
rect 44132 12506 44396 12516
rect 45612 12460 46004 12516
rect 44380 12404 44436 12414
rect 44380 12310 44436 12348
rect 45164 12404 45220 12414
rect 45164 12178 45220 12348
rect 45612 12402 45668 12460
rect 45612 12350 45614 12402
rect 45666 12350 45668 12402
rect 45612 12338 45668 12350
rect 47068 12180 47124 12684
rect 47292 12292 47348 13132
rect 47292 12226 47348 12236
rect 45164 12126 45166 12178
rect 45218 12126 45220 12178
rect 45164 12114 45220 12126
rect 47012 12124 47124 12180
rect 47404 12180 47460 15260
rect 47516 15222 47572 15260
rect 48188 15204 48244 15242
rect 48188 15138 48244 15148
rect 48188 14530 48244 14542
rect 48188 14478 48190 14530
rect 48242 14478 48244 14530
rect 47516 14420 47572 14430
rect 47516 14326 47572 14364
rect 48188 14196 48244 14478
rect 48412 14532 48468 15932
rect 48972 15314 49028 16044
rect 49308 16098 49364 16110
rect 49308 16046 49310 16098
rect 49362 16046 49364 16098
rect 49308 15988 49364 16046
rect 49308 15922 49364 15932
rect 48972 15262 48974 15314
rect 49026 15262 49028 15314
rect 48972 15250 49028 15262
rect 49196 15314 49252 15326
rect 49196 15262 49198 15314
rect 49250 15262 49252 15314
rect 48748 15202 48804 15214
rect 48748 15150 48750 15202
rect 48802 15150 48804 15202
rect 48748 15148 48804 15150
rect 49196 15204 49252 15262
rect 48748 15092 49028 15148
rect 49196 15138 49252 15148
rect 48412 14476 48916 14532
rect 48188 14130 48244 14140
rect 48524 14306 48580 14318
rect 48524 14254 48526 14306
rect 48578 14254 48580 14306
rect 47852 13748 47908 13758
rect 47908 13692 48020 13748
rect 47852 13682 47908 13692
rect 47628 13076 47684 13086
rect 47628 13074 47796 13076
rect 47628 13022 47630 13074
rect 47682 13022 47796 13074
rect 47628 13020 47796 13022
rect 47628 13010 47684 13020
rect 47516 12740 47572 12750
rect 47516 12646 47572 12684
rect 47516 12404 47572 12414
rect 47516 12310 47572 12348
rect 47740 12290 47796 13020
rect 47852 12404 47908 12414
rect 47964 12404 48020 13692
rect 48524 13188 48580 14254
rect 48748 14196 48804 14206
rect 48748 13748 48804 14140
rect 48860 13858 48916 14476
rect 48860 13806 48862 13858
rect 48914 13806 48916 13858
rect 48860 13794 48916 13806
rect 48524 13122 48580 13132
rect 48636 13746 48804 13748
rect 48636 13694 48750 13746
rect 48802 13694 48804 13746
rect 48636 13692 48804 13694
rect 48076 12964 48132 12974
rect 48076 12628 48132 12908
rect 48524 12964 48580 12974
rect 48636 12964 48692 13692
rect 48748 13682 48804 13692
rect 48748 13524 48804 13534
rect 48748 13186 48804 13468
rect 48748 13134 48750 13186
rect 48802 13134 48804 13186
rect 48748 13122 48804 13134
rect 48972 13188 49028 15092
rect 49868 15092 49924 15102
rect 49196 14532 49252 14542
rect 49196 14530 49476 14532
rect 49196 14478 49198 14530
rect 49250 14478 49476 14530
rect 49196 14476 49476 14478
rect 49196 14466 49252 14476
rect 49084 14418 49140 14430
rect 49084 14366 49086 14418
rect 49138 14366 49140 14418
rect 49084 13748 49140 14366
rect 49420 14084 49476 14476
rect 49868 14308 49924 15036
rect 49980 14532 50036 24556
rect 50092 20132 50148 20142
rect 50092 20038 50148 20076
rect 50204 19908 50260 25230
rect 50092 19852 50260 19908
rect 50092 15092 50148 19852
rect 50316 15148 50372 26012
rect 50428 25618 50484 26012
rect 50428 25566 50430 25618
rect 50482 25566 50484 25618
rect 50428 25554 50484 25566
rect 50652 26292 50708 26350
rect 51324 26292 51380 26302
rect 50652 26290 51380 26292
rect 50652 26238 51326 26290
rect 51378 26238 51380 26290
rect 50652 26236 51380 26238
rect 50652 24724 50708 26236
rect 51324 26226 51380 26236
rect 56924 26290 56980 26302
rect 56924 26238 56926 26290
rect 56978 26238 56980 26290
rect 51772 26180 51828 26190
rect 53004 26180 53060 26190
rect 51212 26068 51268 26106
rect 51772 26086 51828 26124
rect 52892 26178 53060 26180
rect 52892 26126 53006 26178
rect 53058 26126 53060 26178
rect 52892 26124 53060 26126
rect 51212 26002 51268 26012
rect 51286 25900 51550 25910
rect 51342 25844 51390 25900
rect 51446 25844 51494 25900
rect 51286 25834 51550 25844
rect 51884 25506 51940 25518
rect 51884 25454 51886 25506
rect 51938 25454 51940 25506
rect 51548 25284 51604 25294
rect 51548 25282 51716 25284
rect 51548 25230 51550 25282
rect 51602 25230 51716 25282
rect 51548 25228 51716 25230
rect 51548 25218 51604 25228
rect 50876 24724 50932 24734
rect 50652 24722 50932 24724
rect 50652 24670 50878 24722
rect 50930 24670 50932 24722
rect 50652 24668 50932 24670
rect 50876 24658 50932 24668
rect 50540 24612 50596 24622
rect 50540 23266 50596 24556
rect 51286 24332 51550 24342
rect 51342 24276 51390 24332
rect 51446 24276 51494 24332
rect 51286 24266 51550 24276
rect 50540 23214 50542 23266
rect 50594 23214 50596 23266
rect 50540 23202 50596 23214
rect 51100 24050 51156 24062
rect 51100 23998 51102 24050
rect 51154 23998 51156 24050
rect 50428 22708 50484 22718
rect 50428 18228 50484 22652
rect 50652 22370 50708 22382
rect 50652 22318 50654 22370
rect 50706 22318 50708 22370
rect 50652 21476 50708 22318
rect 51100 21812 51156 23998
rect 51548 23940 51604 23950
rect 51660 23940 51716 25228
rect 51884 24836 51940 25454
rect 52108 25506 52164 25518
rect 52108 25454 52110 25506
rect 52162 25454 52164 25506
rect 52108 24948 52164 25454
rect 52892 25282 52948 26124
rect 53004 26114 53060 26124
rect 53228 26178 53284 26190
rect 53228 26126 53230 26178
rect 53282 26126 53284 26178
rect 52892 25230 52894 25282
rect 52946 25230 52948 25282
rect 52108 24892 52612 24948
rect 51884 24780 52276 24836
rect 52220 24724 52276 24780
rect 52444 24724 52500 24734
rect 52220 24722 52500 24724
rect 52220 24670 52446 24722
rect 52498 24670 52500 24722
rect 52220 24668 52500 24670
rect 52108 24612 52164 24622
rect 52108 24610 52388 24612
rect 52108 24558 52110 24610
rect 52162 24558 52388 24610
rect 52108 24556 52388 24558
rect 52108 24546 52164 24556
rect 51548 23938 51716 23940
rect 51548 23886 51550 23938
rect 51602 23886 51716 23938
rect 51548 23884 51716 23886
rect 51548 23874 51604 23884
rect 51324 23828 51380 23838
rect 51324 23734 51380 23772
rect 51286 22764 51550 22774
rect 51342 22708 51390 22764
rect 51446 22708 51494 22764
rect 51286 22698 51550 22708
rect 51660 22596 51716 23884
rect 51324 22594 51716 22596
rect 51324 22542 51662 22594
rect 51714 22542 51716 22594
rect 51324 22540 51716 22542
rect 51212 21812 51268 21822
rect 51100 21756 51212 21812
rect 51212 21746 51268 21756
rect 50988 21588 51044 21598
rect 51324 21588 51380 22540
rect 51660 22530 51716 22540
rect 51884 23828 51940 23838
rect 51884 23154 51940 23772
rect 52108 23716 52164 23726
rect 52220 23716 52276 23726
rect 52108 23714 52220 23716
rect 52108 23662 52110 23714
rect 52162 23662 52220 23714
rect 52108 23660 52220 23662
rect 52108 23650 52164 23660
rect 52108 23268 52164 23278
rect 52108 23174 52164 23212
rect 51884 23102 51886 23154
rect 51938 23102 51940 23154
rect 51436 22372 51492 22382
rect 51884 22372 51940 23102
rect 51436 22370 51940 22372
rect 51436 22318 51438 22370
rect 51490 22318 51940 22370
rect 51436 22316 51940 22318
rect 51436 22306 51492 22316
rect 51996 22148 52052 22158
rect 51772 22146 52052 22148
rect 51772 22094 51998 22146
rect 52050 22094 52052 22146
rect 51772 22092 52052 22094
rect 50988 21586 51380 21588
rect 50988 21534 50990 21586
rect 51042 21534 51380 21586
rect 50988 21532 51380 21534
rect 51436 21698 51492 21710
rect 51436 21646 51438 21698
rect 51490 21646 51492 21698
rect 50988 21522 51044 21532
rect 50652 21474 50820 21476
rect 50652 21422 50654 21474
rect 50706 21422 50820 21474
rect 50652 21420 50820 21422
rect 50652 21410 50708 21420
rect 50652 20916 50708 20926
rect 50540 19012 50596 19022
rect 50540 18450 50596 18956
rect 50540 18398 50542 18450
rect 50594 18398 50596 18450
rect 50540 18386 50596 18398
rect 50428 18172 50596 18228
rect 50428 16772 50484 16782
rect 50428 15540 50484 16716
rect 50428 15474 50484 15484
rect 50092 15026 50148 15036
rect 50204 15092 50372 15148
rect 50428 15204 50484 15214
rect 49980 14476 50148 14532
rect 49980 14308 50036 14318
rect 49308 13972 49364 13982
rect 49084 13682 49140 13692
rect 49196 13970 49364 13972
rect 49196 13918 49310 13970
rect 49362 13918 49364 13970
rect 49196 13916 49364 13918
rect 49084 13188 49140 13198
rect 48972 13186 49140 13188
rect 48972 13134 49086 13186
rect 49138 13134 49140 13186
rect 48972 13132 49140 13134
rect 49084 13122 49140 13132
rect 48972 12964 49028 12974
rect 48636 12962 49028 12964
rect 48636 12910 48974 12962
rect 49026 12910 49028 12962
rect 48636 12908 49028 12910
rect 48524 12870 48580 12908
rect 48972 12898 49028 12908
rect 48636 12740 48692 12750
rect 48636 12738 48916 12740
rect 48636 12686 48638 12738
rect 48690 12686 48916 12738
rect 48636 12684 48916 12686
rect 48636 12674 48692 12684
rect 48076 12572 48244 12628
rect 48076 12404 48132 12414
rect 47964 12402 48132 12404
rect 47964 12350 48078 12402
rect 48130 12350 48132 12402
rect 47964 12348 48132 12350
rect 47852 12310 47908 12348
rect 48076 12338 48132 12348
rect 47740 12238 47742 12290
rect 47794 12238 47796 12290
rect 47740 12226 47796 12238
rect 47404 12124 47684 12180
rect 47012 12078 47068 12124
rect 44716 12068 44772 12078
rect 45500 12068 45556 12078
rect 44716 12066 44884 12068
rect 44716 12014 44718 12066
rect 44770 12014 44884 12066
rect 44716 12012 44884 12014
rect 44716 12002 44772 12012
rect 44716 11844 44772 11854
rect 44716 11394 44772 11788
rect 44828 11508 44884 12012
rect 44940 11956 44996 11966
rect 44940 11954 45108 11956
rect 44940 11902 44942 11954
rect 44994 11902 45108 11954
rect 44940 11900 45108 11902
rect 44940 11890 44996 11900
rect 44940 11508 44996 11518
rect 44828 11506 44996 11508
rect 44828 11454 44942 11506
rect 44994 11454 44996 11506
rect 44828 11452 44996 11454
rect 44940 11442 44996 11452
rect 44716 11342 44718 11394
rect 44770 11342 44772 11394
rect 44716 11330 44772 11342
rect 43932 11218 43988 11228
rect 44268 11284 44324 11294
rect 44268 11190 44324 11228
rect 45052 11284 45108 11900
rect 45276 11394 45332 11406
rect 45276 11342 45278 11394
rect 45330 11342 45332 11394
rect 45052 11218 45108 11228
rect 45164 11282 45220 11294
rect 45164 11230 45166 11282
rect 45218 11230 45220 11282
rect 43596 11172 43652 11182
rect 43036 10518 43092 10556
rect 43484 10610 43540 10622
rect 43484 10558 43486 10610
rect 43538 10558 43540 10610
rect 42924 10108 43428 10164
rect 42924 9940 42980 9950
rect 43372 9940 43428 10108
rect 42924 9938 43316 9940
rect 42924 9886 42926 9938
rect 42978 9886 43316 9938
rect 42924 9884 43316 9886
rect 42924 9874 42980 9884
rect 42588 9828 42644 9838
rect 42476 9826 42644 9828
rect 42476 9774 42590 9826
rect 42642 9774 42644 9826
rect 42476 9772 42644 9774
rect 42588 9762 42644 9772
rect 42364 9716 42420 9726
rect 42364 9622 42420 9660
rect 42812 9602 42868 9614
rect 42812 9550 42814 9602
rect 42866 9550 42868 9602
rect 42252 9324 42756 9380
rect 42588 9156 42644 9166
rect 42588 9062 42644 9100
rect 42140 8318 42142 8370
rect 42194 8318 42196 8370
rect 42140 8306 42196 8318
rect 42252 8372 42308 8382
rect 42252 8148 42308 8316
rect 42476 8260 42532 8270
rect 42476 8166 42532 8204
rect 42700 8258 42756 9324
rect 42812 9268 42868 9550
rect 42812 9202 42868 9212
rect 42924 9602 42980 9614
rect 42924 9550 42926 9602
rect 42978 9550 42980 9602
rect 42700 8206 42702 8258
rect 42754 8206 42756 8258
rect 42700 8194 42756 8206
rect 42812 9044 42868 9054
rect 42028 8092 42196 8148
rect 42140 7812 42196 8092
rect 42252 8146 42420 8148
rect 42252 8094 42254 8146
rect 42306 8094 42420 8146
rect 42252 8092 42420 8094
rect 42252 8082 42308 8092
rect 42140 7756 42308 7812
rect 41244 7588 41300 7598
rect 41244 7494 41300 7532
rect 42140 7588 42196 7598
rect 42140 7494 42196 7532
rect 41132 7410 41188 7420
rect 42028 7476 42084 7486
rect 42028 7382 42084 7420
rect 40908 6692 40964 6702
rect 40796 6690 40964 6692
rect 40796 6638 40910 6690
rect 40962 6638 40964 6690
rect 40796 6636 40964 6638
rect 40908 6626 40964 6636
rect 41244 6690 41300 6702
rect 41244 6638 41246 6690
rect 41298 6638 41300 6690
rect 40236 6178 40292 6188
rect 40124 6078 40126 6130
rect 40178 6078 40180 6130
rect 40124 6066 40180 6078
rect 39452 5030 39508 5068
rect 39788 5628 39956 5684
rect 41244 5908 41300 6638
rect 42028 6692 42084 6702
rect 42028 6598 42084 6636
rect 42252 6692 42308 7756
rect 42252 6626 42308 6636
rect 42364 6580 42420 8092
rect 42812 8036 42868 8988
rect 42700 7980 42868 8036
rect 42924 8596 42980 9550
rect 43036 9044 43092 9054
rect 43036 8950 43092 8988
rect 42924 8540 43204 8596
rect 42700 6802 42756 7980
rect 42700 6750 42702 6802
rect 42754 6750 42756 6802
rect 42700 6738 42756 6750
rect 42812 6690 42868 6702
rect 42812 6638 42814 6690
rect 42866 6638 42868 6690
rect 42812 6580 42868 6638
rect 42364 6524 42868 6580
rect 42924 6468 42980 8540
rect 43148 8482 43204 8540
rect 43148 8430 43150 8482
rect 43202 8430 43204 8482
rect 43148 8418 43204 8430
rect 43260 7588 43316 9884
rect 43372 9156 43428 9884
rect 43484 9828 43540 10558
rect 43484 9762 43540 9772
rect 43484 9604 43540 9614
rect 43596 9604 43652 11116
rect 44132 11004 44396 11014
rect 44188 10948 44236 11004
rect 44292 10948 44340 11004
rect 44132 10938 44396 10948
rect 43484 9602 43652 9604
rect 43484 9550 43486 9602
rect 43538 9550 43652 9602
rect 43484 9548 43652 9550
rect 45052 10610 45108 10622
rect 45052 10558 45054 10610
rect 45106 10558 45108 10610
rect 45052 9826 45108 10558
rect 45164 9940 45220 11230
rect 45276 11172 45332 11342
rect 45276 11106 45332 11116
rect 45164 9874 45220 9884
rect 45276 10498 45332 10510
rect 45276 10446 45278 10498
rect 45330 10446 45332 10498
rect 45052 9774 45054 9826
rect 45106 9774 45108 9826
rect 43484 9380 43540 9548
rect 45052 9492 45108 9774
rect 45276 9716 45332 10446
rect 44132 9436 44396 9446
rect 44188 9380 44236 9436
rect 44292 9380 44340 9436
rect 44132 9370 44396 9380
rect 44604 9436 45108 9492
rect 45164 9660 45276 9716
rect 43484 9314 43540 9324
rect 43596 9156 43652 9166
rect 43372 9154 43652 9156
rect 43372 9102 43598 9154
rect 43650 9102 43652 9154
rect 43372 9100 43652 9102
rect 43596 9090 43652 9100
rect 44604 9154 44660 9436
rect 44604 9102 44606 9154
rect 44658 9102 44660 9154
rect 44604 8932 44660 9102
rect 44716 9268 44772 9278
rect 45164 9268 45220 9660
rect 45276 9650 45332 9660
rect 44716 9042 44772 9212
rect 44716 8990 44718 9042
rect 44770 8990 44772 9042
rect 44716 8978 44772 8990
rect 45052 9212 45220 9268
rect 45388 9380 45444 9390
rect 44604 8866 44660 8876
rect 43484 8260 43540 8270
rect 45052 8260 45108 9212
rect 45276 9156 45332 9166
rect 43484 8166 43540 8204
rect 44940 8258 45108 8260
rect 44940 8206 45054 8258
rect 45106 8206 45108 8258
rect 44940 8204 45108 8206
rect 43260 7522 43316 7532
rect 43372 8146 43428 8158
rect 43372 8094 43374 8146
rect 43426 8094 43428 8146
rect 43148 6916 43204 6926
rect 43148 6822 43204 6860
rect 42140 6412 42980 6468
rect 43036 6692 43092 6702
rect 42140 6130 42196 6412
rect 42140 6078 42142 6130
rect 42194 6078 42196 6130
rect 42140 6066 42196 6078
rect 39788 5122 39844 5628
rect 40348 5460 40404 5470
rect 39788 5070 39790 5122
rect 39842 5070 39844 5122
rect 39788 5058 39844 5070
rect 40012 5124 40068 5134
rect 39900 5010 39956 5022
rect 39900 4958 39902 5010
rect 39954 4958 39956 5010
rect 39900 4900 39956 4958
rect 39228 4844 39956 4900
rect 40012 4898 40068 5068
rect 40012 4846 40014 4898
rect 40066 4846 40068 4898
rect 39228 4338 39284 4844
rect 40012 4834 40068 4846
rect 40348 4562 40404 5404
rect 40684 5124 40740 5134
rect 40684 5030 40740 5068
rect 40348 4510 40350 4562
rect 40402 4510 40404 4562
rect 40348 4452 40404 4510
rect 40348 4386 40404 4396
rect 41244 4340 41300 5852
rect 42028 5906 42084 5918
rect 42028 5854 42030 5906
rect 42082 5854 42084 5906
rect 41580 5236 41636 5246
rect 42028 5236 42084 5854
rect 41580 5142 41636 5180
rect 41916 5180 42084 5236
rect 41916 4900 41972 5180
rect 42140 5124 42196 5134
rect 39228 4286 39230 4338
rect 39282 4286 39284 4338
rect 39228 4274 39284 4286
rect 41132 4338 41300 4340
rect 41132 4286 41246 4338
rect 41298 4286 41300 4338
rect 41132 4284 41300 4286
rect 39004 4174 39006 4226
rect 39058 4174 39060 4226
rect 39004 4162 39060 4174
rect 38108 3490 38164 3500
rect 41132 3556 41188 4284
rect 41244 4274 41300 4284
rect 41356 4452 41412 4462
rect 41244 3668 41300 3678
rect 41356 3668 41412 4396
rect 41580 4340 41636 4350
rect 41580 4246 41636 4284
rect 41244 3666 41356 3668
rect 41244 3614 41246 3666
rect 41298 3614 41356 3666
rect 41244 3612 41356 3614
rect 41244 3602 41300 3612
rect 41356 3574 41412 3612
rect 41132 3490 41188 3500
rect 41468 3556 41524 3566
rect 41468 3462 41524 3500
rect 37660 3442 38052 3444
rect 37660 3390 37662 3442
rect 37714 3390 38052 3442
rect 37660 3388 38052 3390
rect 41916 3442 41972 4844
rect 42028 5068 42140 5124
rect 42028 3666 42084 5068
rect 42140 5058 42196 5068
rect 42028 3614 42030 3666
rect 42082 3614 42084 3666
rect 42028 3602 42084 3614
rect 42364 3668 42420 3678
rect 42364 3554 42420 3612
rect 42364 3502 42366 3554
rect 42418 3502 42420 3554
rect 42364 3490 42420 3502
rect 41916 3390 41918 3442
rect 41970 3390 41972 3442
rect 37660 3378 37716 3388
rect 41916 3378 41972 3390
rect 42476 3444 42532 6412
rect 43036 6132 43092 6636
rect 43036 6018 43092 6076
rect 43036 5966 43038 6018
rect 43090 5966 43092 6018
rect 43036 5954 43092 5966
rect 42812 5908 42868 5918
rect 42812 5814 42868 5852
rect 42700 5794 42756 5806
rect 42700 5742 42702 5794
rect 42754 5742 42756 5794
rect 42588 4340 42644 4350
rect 42700 4340 42756 5742
rect 43372 5234 43428 8094
rect 44044 8148 44100 8158
rect 44828 8148 44884 8158
rect 44044 8146 44884 8148
rect 44044 8094 44046 8146
rect 44098 8094 44830 8146
rect 44882 8094 44884 8146
rect 44044 8092 44884 8094
rect 44044 8082 44100 8092
rect 44132 7868 44396 7878
rect 44188 7812 44236 7868
rect 44292 7812 44340 7868
rect 44132 7802 44396 7812
rect 43596 7698 43652 7710
rect 43596 7646 43598 7698
rect 43650 7646 43652 7698
rect 43596 6468 43652 7646
rect 44716 7586 44772 8092
rect 44828 8082 44884 8092
rect 44716 7534 44718 7586
rect 44770 7534 44772 7586
rect 44716 7522 44772 7534
rect 43708 7474 43764 7486
rect 43708 7422 43710 7474
rect 43762 7422 43764 7474
rect 43708 6804 43764 7422
rect 44268 7476 44324 7486
rect 43932 6916 43988 6926
rect 43932 6822 43988 6860
rect 44268 6914 44324 7420
rect 44940 7252 44996 8204
rect 45052 8194 45108 8204
rect 45164 9100 45276 9156
rect 45164 8146 45220 9100
rect 45276 9090 45332 9100
rect 45388 8260 45444 9324
rect 45500 8820 45556 12012
rect 46956 12066 47068 12078
rect 46956 12014 46958 12066
rect 47010 12014 47068 12066
rect 46956 12012 47068 12014
rect 46956 11844 47012 12012
rect 46620 11788 47012 11844
rect 45948 11508 46004 11518
rect 46004 11452 46452 11508
rect 45948 11414 46004 11452
rect 46284 11170 46340 11182
rect 46284 11118 46286 11170
rect 46338 11118 46340 11170
rect 46284 10500 46340 11118
rect 46396 10724 46452 11452
rect 46396 10630 46452 10668
rect 46620 10722 46676 11788
rect 47516 11732 47572 11742
rect 47516 11508 47572 11676
rect 46956 11506 47572 11508
rect 46956 11454 47518 11506
rect 47570 11454 47572 11506
rect 46956 11452 47572 11454
rect 46844 11284 46900 11294
rect 46620 10670 46622 10722
rect 46674 10670 46676 10722
rect 46284 10434 46340 10444
rect 46620 10500 46676 10670
rect 46620 10434 46676 10444
rect 46732 11282 46900 11284
rect 46732 11230 46846 11282
rect 46898 11230 46900 11282
rect 46732 11228 46900 11230
rect 46732 10498 46788 11228
rect 46844 11218 46900 11228
rect 46956 11282 47012 11452
rect 46956 11230 46958 11282
rect 47010 11230 47012 11282
rect 46956 11218 47012 11230
rect 47068 11284 47124 11294
rect 47124 11228 47236 11284
rect 47068 11218 47124 11228
rect 47180 11170 47236 11228
rect 47180 11118 47182 11170
rect 47234 11118 47236 11170
rect 47180 11106 47236 11118
rect 47292 10722 47348 11452
rect 47516 11442 47572 11452
rect 47628 10724 47684 12124
rect 48188 11508 48244 12572
rect 48524 12516 48580 12526
rect 47964 11452 48244 11508
rect 48300 12292 48356 12302
rect 48300 11956 48356 12236
rect 48300 11506 48356 11900
rect 48300 11454 48302 11506
rect 48354 11454 48356 11506
rect 47964 11172 48020 11452
rect 48300 11442 48356 11454
rect 48076 11284 48132 11294
rect 48132 11228 48244 11284
rect 48076 11218 48132 11228
rect 47292 10670 47294 10722
rect 47346 10670 47348 10722
rect 47292 10658 47348 10670
rect 47516 10668 47684 10724
rect 47852 10724 47908 10734
rect 47404 10610 47460 10622
rect 47404 10558 47406 10610
rect 47458 10558 47460 10610
rect 46732 10446 46734 10498
rect 46786 10446 46788 10498
rect 46732 10434 46788 10446
rect 47068 10500 47124 10510
rect 46956 9940 47012 9950
rect 46956 9846 47012 9884
rect 46732 9826 46788 9838
rect 46732 9774 46734 9826
rect 46786 9774 46788 9826
rect 46508 9716 46564 9726
rect 46508 9622 46564 9660
rect 46396 9156 46452 9166
rect 46732 9156 46788 9774
rect 47068 9266 47124 10444
rect 47404 10500 47460 10558
rect 47404 10434 47460 10444
rect 47068 9214 47070 9266
rect 47122 9214 47124 9266
rect 47068 9202 47124 9214
rect 46396 9154 46732 9156
rect 46396 9102 46398 9154
rect 46450 9102 46732 9154
rect 46396 9100 46732 9102
rect 46396 9090 46452 9100
rect 46732 9090 46788 9100
rect 47516 9044 47572 10668
rect 47852 10610 47908 10668
rect 47852 10558 47854 10610
rect 47906 10558 47908 10610
rect 47852 10546 47908 10558
rect 47628 10498 47684 10510
rect 47628 10446 47630 10498
rect 47682 10446 47684 10498
rect 47628 9828 47684 10446
rect 47964 10052 48020 11116
rect 47964 9958 48020 9996
rect 48076 10386 48132 10398
rect 48076 10334 48078 10386
rect 48130 10334 48132 10386
rect 47628 9762 47684 9772
rect 47068 8988 47572 9044
rect 47628 9604 47684 9614
rect 47628 9044 47684 9548
rect 48076 9602 48132 10334
rect 48188 10052 48244 11228
rect 48524 10052 48580 12460
rect 48636 12180 48692 12190
rect 48636 11170 48692 12124
rect 48860 12178 48916 12684
rect 49196 12180 49252 13916
rect 49308 13906 49364 13916
rect 49420 13524 49476 14028
rect 49420 13458 49476 13468
rect 49756 14306 50036 14308
rect 49756 14254 49982 14306
rect 50034 14254 50036 14306
rect 49756 14252 50036 14254
rect 49756 12628 49812 14252
rect 49980 14242 50036 14252
rect 49868 14084 49924 14094
rect 49868 13746 49924 14028
rect 49868 13694 49870 13746
rect 49922 13694 49924 13746
rect 49868 13682 49924 13694
rect 50092 13300 50148 14476
rect 49980 13244 50148 13300
rect 49980 13186 50036 13244
rect 50204 13188 50260 15092
rect 50428 14756 50484 15148
rect 50428 14690 50484 14700
rect 50540 14532 50596 18172
rect 50652 15876 50708 20860
rect 50764 20804 50820 21420
rect 51436 21364 51492 21646
rect 51436 21308 51716 21364
rect 51286 21196 51550 21206
rect 51342 21140 51390 21196
rect 51446 21140 51494 21196
rect 51286 21130 51550 21140
rect 50764 17668 50820 20748
rect 51548 20804 51604 20814
rect 51660 20804 51716 21308
rect 51548 20802 51716 20804
rect 51548 20750 51550 20802
rect 51602 20750 51716 20802
rect 51548 20748 51716 20750
rect 51548 20738 51604 20748
rect 50876 20690 50932 20702
rect 50876 20638 50878 20690
rect 50930 20638 50932 20690
rect 50876 20244 50932 20638
rect 50876 20018 50932 20188
rect 50876 19966 50878 20018
rect 50930 19966 50932 20018
rect 50876 19954 50932 19966
rect 51100 20018 51156 20030
rect 51100 19966 51102 20018
rect 51154 19966 51156 20018
rect 51100 19796 51156 19966
rect 51100 19730 51156 19740
rect 51286 19628 51550 19638
rect 51342 19572 51390 19628
rect 51446 19572 51494 19628
rect 51286 19562 51550 19572
rect 51660 19346 51716 20748
rect 51660 19294 51662 19346
rect 51714 19294 51716 19346
rect 51660 19282 51716 19294
rect 51772 19348 51828 22092
rect 51996 22082 52052 22092
rect 51996 21588 52052 21598
rect 51772 19282 51828 19292
rect 51884 20916 51940 20926
rect 51884 20690 51940 20860
rect 51884 20638 51886 20690
rect 51938 20638 51940 20690
rect 50876 19236 50932 19246
rect 50876 19142 50932 19180
rect 51884 19124 51940 20638
rect 51548 19068 51940 19124
rect 51996 20578 52052 21532
rect 52108 21028 52164 21038
rect 52220 21028 52276 23660
rect 52332 23154 52388 24556
rect 52444 23268 52500 24668
rect 52444 23174 52500 23212
rect 52556 23604 52612 24892
rect 52892 23828 52948 25230
rect 53004 25508 53060 25518
rect 53228 25508 53284 26126
rect 56588 26180 56644 26190
rect 56924 26180 56980 26238
rect 56588 26178 56980 26180
rect 56588 26126 56590 26178
rect 56642 26126 56980 26178
rect 56588 26124 56980 26126
rect 53452 26068 53508 26078
rect 53452 26066 53620 26068
rect 53452 26014 53454 26066
rect 53506 26014 53620 26066
rect 53452 26012 53620 26014
rect 53452 26002 53508 26012
rect 53564 25618 53620 26012
rect 53564 25566 53566 25618
rect 53618 25566 53620 25618
rect 53452 25508 53508 25518
rect 53228 25506 53508 25508
rect 53228 25454 53454 25506
rect 53506 25454 53508 25506
rect 53228 25452 53508 25454
rect 53004 24834 53060 25452
rect 53004 24782 53006 24834
rect 53058 24782 53060 24834
rect 53004 24770 53060 24782
rect 52892 23762 52948 23772
rect 53116 23940 53172 23950
rect 53340 23940 53396 25452
rect 53452 25442 53508 25452
rect 53116 23938 53396 23940
rect 53116 23886 53118 23938
rect 53170 23886 53396 23938
rect 53116 23884 53396 23886
rect 53452 24610 53508 24622
rect 53452 24558 53454 24610
rect 53506 24558 53508 24610
rect 53116 23604 53172 23884
rect 52556 23548 53172 23604
rect 52332 23102 52334 23154
rect 52386 23102 52388 23154
rect 52332 22932 52388 23102
rect 52332 22866 52388 22876
rect 52164 20972 52276 21028
rect 52332 21810 52388 21822
rect 52332 21758 52334 21810
rect 52386 21758 52388 21810
rect 52108 20962 52164 20972
rect 52220 20692 52276 20702
rect 52220 20598 52276 20636
rect 51996 20526 51998 20578
rect 52050 20526 52052 20578
rect 51548 18788 51604 19068
rect 51548 18732 51828 18788
rect 51286 18060 51550 18070
rect 51342 18004 51390 18060
rect 51446 18004 51494 18060
rect 51286 17994 51550 18004
rect 50876 17668 50932 17678
rect 50764 17666 50932 17668
rect 50764 17614 50878 17666
rect 50930 17614 50932 17666
rect 50764 17612 50932 17614
rect 50876 17602 50932 17612
rect 51212 17444 51268 17454
rect 51660 17444 51716 17454
rect 51212 17442 51380 17444
rect 51212 17390 51214 17442
rect 51266 17390 51380 17442
rect 51212 17388 51380 17390
rect 51212 17378 51268 17388
rect 50652 15810 50708 15820
rect 50988 16996 51044 17006
rect 50652 15428 50708 15438
rect 50988 15428 51044 16940
rect 51324 16882 51380 17388
rect 51324 16830 51326 16882
rect 51378 16830 51380 16882
rect 51324 16660 51380 16830
rect 51548 17388 51660 17444
rect 51548 16772 51604 17388
rect 51660 17350 51716 17388
rect 51772 17220 51828 18732
rect 51548 16706 51604 16716
rect 51660 17164 51828 17220
rect 51884 18674 51940 18686
rect 51884 18622 51886 18674
rect 51938 18622 51940 18674
rect 51100 16604 51380 16660
rect 51100 16098 51156 16604
rect 51286 16492 51550 16502
rect 51342 16436 51390 16492
rect 51446 16436 51494 16492
rect 51286 16426 51550 16436
rect 51660 16324 51716 17164
rect 51884 16994 51940 18622
rect 51996 17444 52052 20526
rect 52332 18564 52388 21758
rect 52444 19796 52500 19806
rect 52556 19796 52612 23548
rect 53452 23492 53508 24558
rect 53564 23938 53620 25566
rect 53676 26066 53732 26078
rect 53676 26014 53678 26066
rect 53730 26014 53732 26066
rect 53676 25508 53732 26014
rect 53676 25442 53732 25452
rect 54124 26066 54180 26078
rect 54124 26014 54126 26066
rect 54178 26014 54180 26066
rect 54124 24724 54180 26014
rect 54908 25730 54964 25742
rect 54908 25678 54910 25730
rect 54962 25678 54964 25730
rect 54908 24834 54964 25678
rect 56588 25620 56644 26124
rect 56588 25554 56644 25564
rect 55468 25508 55524 25518
rect 55468 25414 55524 25452
rect 58439 25116 58703 25126
rect 58495 25060 58543 25116
rect 58599 25060 58647 25116
rect 58439 25050 58703 25060
rect 54908 24782 54910 24834
rect 54962 24782 54964 24834
rect 54572 24724 54628 24734
rect 54124 24722 54628 24724
rect 54124 24670 54574 24722
rect 54626 24670 54628 24722
rect 54124 24668 54628 24670
rect 54572 24658 54628 24668
rect 53564 23886 53566 23938
rect 53618 23886 53620 23938
rect 53564 23716 53620 23886
rect 54908 23940 54964 24782
rect 55244 24612 55300 24622
rect 55244 24610 55412 24612
rect 55244 24558 55246 24610
rect 55298 24558 55412 24610
rect 55244 24556 55412 24558
rect 55244 24546 55300 24556
rect 54908 23874 54964 23884
rect 54236 23828 54292 23838
rect 53564 23650 53620 23660
rect 54012 23826 54292 23828
rect 54012 23774 54238 23826
rect 54290 23774 54292 23826
rect 54012 23772 54292 23774
rect 53116 23436 53508 23492
rect 52668 23380 52724 23390
rect 52668 23286 52724 23324
rect 53004 23044 53060 23054
rect 53116 23044 53172 23436
rect 53004 23042 53172 23044
rect 53004 22990 53006 23042
rect 53058 22990 53172 23042
rect 53004 22988 53172 22990
rect 53228 23268 53284 23278
rect 53004 22932 53060 22988
rect 53004 22866 53060 22876
rect 52780 22596 52836 22606
rect 52780 22370 52836 22540
rect 52780 22318 52782 22370
rect 52834 22318 52836 22370
rect 52780 21812 52836 22318
rect 53004 22484 53060 22494
rect 53004 22370 53060 22428
rect 53004 22318 53006 22370
rect 53058 22318 53060 22370
rect 52892 22148 52948 22158
rect 52892 22054 52948 22092
rect 52780 21756 52948 21812
rect 52780 21474 52836 21486
rect 52780 21422 52782 21474
rect 52834 21422 52836 21474
rect 52668 20802 52724 20814
rect 52668 20750 52670 20802
rect 52722 20750 52724 20802
rect 52668 20468 52724 20750
rect 52668 20402 52724 20412
rect 52780 20020 52836 21422
rect 52892 20914 52948 21756
rect 52892 20862 52894 20914
rect 52946 20862 52948 20914
rect 52892 20850 52948 20862
rect 53004 20804 53060 22318
rect 53228 22258 53284 23212
rect 53452 23154 53508 23166
rect 53452 23102 53454 23154
rect 53506 23102 53508 23154
rect 53228 22206 53230 22258
rect 53282 22206 53284 22258
rect 53228 22194 53284 22206
rect 53340 22372 53396 22382
rect 53340 21924 53396 22316
rect 53452 22260 53508 23102
rect 53676 23156 53732 23166
rect 54012 23156 54068 23772
rect 54236 23762 54292 23772
rect 54796 23716 54852 23726
rect 54684 23714 54852 23716
rect 54684 23662 54798 23714
rect 54850 23662 54852 23714
rect 54684 23660 54852 23662
rect 54572 23604 54628 23614
rect 53676 23154 54068 23156
rect 53676 23102 53678 23154
rect 53730 23102 54068 23154
rect 53676 23100 54068 23102
rect 54124 23154 54180 23166
rect 54124 23102 54126 23154
rect 54178 23102 54180 23154
rect 53676 23090 53732 23100
rect 53452 22194 53508 22204
rect 53564 23042 53620 23054
rect 53564 22990 53566 23042
rect 53618 22990 53620 23042
rect 53340 21868 53508 21924
rect 53340 21586 53396 21598
rect 53340 21534 53342 21586
rect 53394 21534 53396 21586
rect 53116 20804 53172 20814
rect 53004 20802 53172 20804
rect 53004 20750 53118 20802
rect 53170 20750 53172 20802
rect 53004 20748 53172 20750
rect 52780 19954 52836 19964
rect 52892 20244 52948 20254
rect 52892 20018 52948 20188
rect 52892 19966 52894 20018
rect 52946 19966 52948 20018
rect 52500 19740 52612 19796
rect 52444 19730 52500 19740
rect 52332 18470 52388 18508
rect 52556 18452 52612 18462
rect 52556 18358 52612 18396
rect 52892 17780 52948 19966
rect 53004 19236 53060 20748
rect 53116 20738 53172 20748
rect 53228 20580 53284 20590
rect 53228 20486 53284 20524
rect 53340 20578 53396 21534
rect 53452 21252 53508 21868
rect 53564 21700 53620 22990
rect 53788 22372 53844 23100
rect 53564 21634 53620 21644
rect 53676 22260 53732 22270
rect 53676 21364 53732 22204
rect 53788 22258 53844 22316
rect 53788 22206 53790 22258
rect 53842 22206 53844 22258
rect 53788 22194 53844 22206
rect 54012 22146 54068 22158
rect 54012 22094 54014 22146
rect 54066 22094 54068 22146
rect 54012 21924 54068 22094
rect 53788 21868 54068 21924
rect 53788 21586 53844 21868
rect 54124 21812 54180 23102
rect 54348 22370 54404 22382
rect 54348 22318 54350 22370
rect 54402 22318 54404 22370
rect 54348 22260 54404 22318
rect 54348 22194 54404 22204
rect 54124 21746 54180 21756
rect 54236 21810 54292 21822
rect 54236 21758 54238 21810
rect 54290 21758 54292 21810
rect 53788 21534 53790 21586
rect 53842 21534 53844 21586
rect 53788 21522 53844 21534
rect 53900 21698 53956 21710
rect 53900 21646 53902 21698
rect 53954 21646 53956 21698
rect 53900 21588 53956 21646
rect 53900 21522 53956 21532
rect 53676 21308 53956 21364
rect 53452 21196 53844 21252
rect 53788 20914 53844 21196
rect 53788 20862 53790 20914
rect 53842 20862 53844 20914
rect 53788 20850 53844 20862
rect 53340 20526 53342 20578
rect 53394 20526 53396 20578
rect 53340 20244 53396 20526
rect 53340 20178 53396 20188
rect 53452 20804 53508 20814
rect 53900 20804 53956 21308
rect 54012 20804 54068 20814
rect 53900 20802 54068 20804
rect 53900 20750 54014 20802
rect 54066 20750 54068 20802
rect 53900 20748 54068 20750
rect 53452 19458 53508 20748
rect 54012 20132 54068 20748
rect 54012 20038 54068 20076
rect 53452 19406 53454 19458
rect 53506 19406 53508 19458
rect 53452 19394 53508 19406
rect 53564 20018 53620 20030
rect 53564 19966 53566 20018
rect 53618 19966 53620 20018
rect 53004 19170 53060 19180
rect 53116 19346 53172 19358
rect 53116 19294 53118 19346
rect 53170 19294 53172 19346
rect 53116 17780 53172 19294
rect 53340 19348 53396 19358
rect 53228 19234 53284 19246
rect 53228 19182 53230 19234
rect 53282 19182 53284 19234
rect 53228 17892 53284 19182
rect 53340 19234 53396 19292
rect 53340 19182 53342 19234
rect 53394 19182 53396 19234
rect 53340 19170 53396 19182
rect 53564 18788 53620 19966
rect 53228 17826 53284 17836
rect 53340 18732 53620 18788
rect 53900 20018 53956 20030
rect 53900 19966 53902 20018
rect 53954 19966 53956 20018
rect 52780 17724 53060 17780
rect 52780 17666 52836 17724
rect 52780 17614 52782 17666
rect 52834 17614 52836 17666
rect 52780 17602 52836 17614
rect 51996 17378 52052 17388
rect 52892 17554 52948 17566
rect 52892 17502 52894 17554
rect 52946 17502 52948 17554
rect 51884 16942 51886 16994
rect 51938 16942 51940 16994
rect 51548 16268 51716 16324
rect 51772 16772 51828 16782
rect 51436 16212 51492 16222
rect 51436 16118 51492 16156
rect 51100 16046 51102 16098
rect 51154 16046 51156 16098
rect 51100 15764 51156 16046
rect 51100 15708 51492 15764
rect 50652 15426 51044 15428
rect 50652 15374 50654 15426
rect 50706 15374 50990 15426
rect 51042 15374 51044 15426
rect 50652 15372 51044 15374
rect 50652 15316 50708 15372
rect 50988 15362 51044 15372
rect 51436 15428 51492 15708
rect 50652 15250 50708 15260
rect 51212 15316 51268 15326
rect 51212 15222 51268 15260
rect 51436 15314 51492 15372
rect 51436 15262 51438 15314
rect 51490 15262 51492 15314
rect 51436 15250 51492 15262
rect 51548 15148 51604 16268
rect 51660 16100 51716 16110
rect 51660 15314 51716 16044
rect 51660 15262 51662 15314
rect 51714 15262 51716 15314
rect 51660 15250 51716 15262
rect 51772 15988 51828 16716
rect 51884 16100 51940 16942
rect 51884 16034 51940 16044
rect 52108 16996 52164 17006
rect 52108 16098 52164 16940
rect 52108 16046 52110 16098
rect 52162 16046 52164 16098
rect 52108 16034 52164 16046
rect 51772 15316 51828 15932
rect 52108 15540 52164 15550
rect 52892 15540 52948 17502
rect 53004 15988 53060 17724
rect 53116 17686 53172 17724
rect 53340 17668 53396 18732
rect 53900 18676 53956 19966
rect 54236 19348 54292 21758
rect 54460 21700 54516 21710
rect 54348 21698 54516 21700
rect 54348 21646 54462 21698
rect 54514 21646 54516 21698
rect 54348 21644 54516 21646
rect 54348 21026 54404 21644
rect 54460 21634 54516 21644
rect 54348 20974 54350 21026
rect 54402 20974 54404 21026
rect 54348 20962 54404 20974
rect 53228 17666 53396 17668
rect 53228 17614 53342 17666
rect 53394 17614 53396 17666
rect 53228 17612 53396 17614
rect 53228 16212 53284 17612
rect 53340 17602 53396 17612
rect 53452 18620 53956 18676
rect 54012 19292 54292 19348
rect 54460 19348 54516 19358
rect 53452 17106 53508 18620
rect 53900 18450 53956 18462
rect 53900 18398 53902 18450
rect 53954 18398 53956 18450
rect 53900 18340 53956 18398
rect 53900 18274 53956 18284
rect 54012 18116 54068 19292
rect 54348 19234 54404 19246
rect 54348 19182 54350 19234
rect 54402 19182 54404 19234
rect 53788 18060 54068 18116
rect 54236 18340 54292 18350
rect 54348 18340 54404 19182
rect 54460 19122 54516 19292
rect 54460 19070 54462 19122
rect 54514 19070 54516 19122
rect 54460 18564 54516 19070
rect 54460 18470 54516 18508
rect 54572 18340 54628 23548
rect 54684 23042 54740 23660
rect 54796 23650 54852 23660
rect 54684 22990 54686 23042
rect 54738 22990 54740 23042
rect 54684 20916 54740 22990
rect 54796 23154 54852 23166
rect 54796 23102 54798 23154
rect 54850 23102 54852 23154
rect 54796 21588 54852 23102
rect 54796 21522 54852 21532
rect 55132 22372 55188 22382
rect 54796 20916 54852 20926
rect 54684 20860 54796 20916
rect 54796 20822 54852 20860
rect 55020 20804 55076 20814
rect 55020 20710 55076 20748
rect 55132 20018 55188 22316
rect 55356 22260 55412 24556
rect 56588 24610 56644 24622
rect 56588 24558 56590 24610
rect 56642 24558 56644 24610
rect 55580 23940 55636 23950
rect 55580 23846 55636 23884
rect 56588 23940 56644 24558
rect 56812 24500 56868 24510
rect 56812 24498 57092 24500
rect 56812 24446 56814 24498
rect 56866 24446 57092 24498
rect 56812 24444 57092 24446
rect 56812 24434 56868 24444
rect 56588 23938 56980 23940
rect 56588 23886 56590 23938
rect 56642 23886 56980 23938
rect 56588 23884 56980 23886
rect 56588 23874 56644 23884
rect 55804 23826 55860 23838
rect 55804 23774 55806 23826
rect 55858 23774 55860 23826
rect 55804 23380 55860 23774
rect 56476 23716 56532 23726
rect 56476 23714 56868 23716
rect 56476 23662 56478 23714
rect 56530 23662 56868 23714
rect 56476 23660 56868 23662
rect 56476 23650 56532 23660
rect 55804 23314 55860 23324
rect 55468 23268 55524 23278
rect 55468 23174 55524 23212
rect 55916 23044 55972 23054
rect 55916 23042 56084 23044
rect 55916 22990 55918 23042
rect 55970 22990 56084 23042
rect 55916 22988 56084 22990
rect 55916 22978 55972 22988
rect 55468 22260 55524 22270
rect 55356 22258 55524 22260
rect 55356 22206 55470 22258
rect 55522 22206 55524 22258
rect 55356 22204 55524 22206
rect 55356 21812 55412 22204
rect 55468 22194 55524 22204
rect 55244 21588 55300 21598
rect 55244 21494 55300 21532
rect 55244 21026 55300 21038
rect 55244 20974 55246 21026
rect 55298 20974 55300 21026
rect 55244 20356 55300 20974
rect 55356 20468 55412 21756
rect 55468 21700 55524 21710
rect 55468 21586 55524 21644
rect 56028 21698 56084 22988
rect 56364 22372 56420 22382
rect 56364 22278 56420 22316
rect 56028 21646 56030 21698
rect 56082 21646 56084 21698
rect 55468 21534 55470 21586
rect 55522 21534 55524 21586
rect 55468 21522 55524 21534
rect 55804 21588 55860 21598
rect 55692 21364 55748 21374
rect 55580 21362 55748 21364
rect 55580 21310 55694 21362
rect 55746 21310 55748 21362
rect 55580 21308 55748 21310
rect 55356 20412 55524 20468
rect 55244 20300 55412 20356
rect 55132 19966 55134 20018
rect 55186 19966 55188 20018
rect 55132 19954 55188 19966
rect 55244 20132 55300 20142
rect 55244 20018 55300 20076
rect 55244 19966 55246 20018
rect 55298 19966 55300 20018
rect 55244 19954 55300 19966
rect 54796 19236 54852 19246
rect 54796 18450 54852 19180
rect 54796 18398 54798 18450
rect 54850 18398 54852 18450
rect 54796 18386 54852 18398
rect 54908 18788 54964 18798
rect 55356 18788 55412 20300
rect 55468 20018 55524 20412
rect 55468 19966 55470 20018
rect 55522 19966 55524 20018
rect 55468 19954 55524 19966
rect 54908 18450 54964 18732
rect 54908 18398 54910 18450
rect 54962 18398 54964 18450
rect 54908 18386 54964 18398
rect 55020 18732 55412 18788
rect 54292 18284 54404 18340
rect 54460 18284 54628 18340
rect 53564 17780 53620 17790
rect 53564 17554 53620 17724
rect 53564 17502 53566 17554
rect 53618 17502 53620 17554
rect 53564 17490 53620 17502
rect 53452 17054 53454 17106
rect 53506 17054 53508 17106
rect 53452 17042 53508 17054
rect 53564 17108 53620 17118
rect 53340 16882 53396 16894
rect 53340 16830 53342 16882
rect 53394 16830 53396 16882
rect 53340 16772 53396 16830
rect 53340 16706 53396 16716
rect 53228 16146 53284 16156
rect 53228 15988 53284 15998
rect 53004 15986 53284 15988
rect 53004 15934 53230 15986
rect 53282 15934 53284 15986
rect 53004 15932 53284 15934
rect 53228 15922 53284 15932
rect 53452 15986 53508 15998
rect 53452 15934 53454 15986
rect 53506 15934 53508 15986
rect 53452 15540 53508 15934
rect 52108 15538 53508 15540
rect 52108 15486 52110 15538
rect 52162 15486 53508 15538
rect 52108 15484 53508 15486
rect 52108 15474 52164 15484
rect 51772 15250 51828 15260
rect 53452 15316 53508 15326
rect 53452 15222 53508 15260
rect 51548 15092 51828 15148
rect 51286 14924 51550 14934
rect 51342 14868 51390 14924
rect 51446 14868 51494 14924
rect 51286 14858 51550 14868
rect 50428 14476 50596 14532
rect 50876 14530 50932 14542
rect 51212 14532 51268 14542
rect 50876 14478 50878 14530
rect 50930 14478 50932 14530
rect 50316 13858 50372 13870
rect 50316 13806 50318 13858
rect 50370 13806 50372 13858
rect 50316 13748 50372 13806
rect 50316 13682 50372 13692
rect 49980 13134 49982 13186
rect 50034 13134 50036 13186
rect 49868 12738 49924 12750
rect 49868 12686 49870 12738
rect 49922 12686 49924 12738
rect 49868 12628 49924 12686
rect 49532 12572 49924 12628
rect 48860 12126 48862 12178
rect 48914 12126 48916 12178
rect 48860 12114 48916 12126
rect 48972 12124 49252 12180
rect 49420 12180 49476 12190
rect 48636 11118 48638 11170
rect 48690 11118 48692 11170
rect 48636 10500 48692 11118
rect 48860 10724 48916 10734
rect 48860 10630 48916 10668
rect 48636 10434 48692 10444
rect 48188 9996 48356 10052
rect 48524 9996 48804 10052
rect 48076 9550 48078 9602
rect 48130 9550 48132 9602
rect 48076 9538 48132 9550
rect 48188 9826 48244 9838
rect 48188 9774 48190 9826
rect 48242 9774 48244 9826
rect 48188 9380 48244 9774
rect 47964 9324 48244 9380
rect 47628 9042 47796 9044
rect 47628 8990 47630 9042
rect 47682 8990 47796 9042
rect 47628 8988 47796 8990
rect 45500 8754 45556 8764
rect 45948 8820 46004 8830
rect 45948 8370 46004 8764
rect 45948 8318 45950 8370
rect 46002 8318 46004 8370
rect 45948 8306 46004 8318
rect 45388 8194 45444 8204
rect 46396 8258 46452 8270
rect 46396 8206 46398 8258
rect 46450 8206 46452 8258
rect 45164 8094 45166 8146
rect 45218 8094 45220 8146
rect 45164 8082 45220 8094
rect 45276 8036 45332 8046
rect 45836 8036 45892 8046
rect 46060 8036 46116 8046
rect 45276 7698 45332 7980
rect 45276 7646 45278 7698
rect 45330 7646 45332 7698
rect 45276 7634 45332 7646
rect 45388 8034 45892 8036
rect 45388 7982 45838 8034
rect 45890 7982 45892 8034
rect 45388 7980 45892 7982
rect 45052 7588 45108 7598
rect 45052 7494 45108 7532
rect 45388 7362 45444 7980
rect 45836 7970 45892 7980
rect 45948 8034 46116 8036
rect 45948 7982 46062 8034
rect 46114 7982 46116 8034
rect 45948 7980 46116 7982
rect 45836 7588 45892 7598
rect 45948 7588 46004 7980
rect 46060 7970 46116 7980
rect 46060 7700 46116 7710
rect 46396 7700 46452 8206
rect 46844 8146 46900 8158
rect 46844 8094 46846 8146
rect 46898 8094 46900 8146
rect 46732 8036 46788 8046
rect 46732 7942 46788 7980
rect 46844 7700 46900 8094
rect 46060 7698 46452 7700
rect 46060 7646 46062 7698
rect 46114 7646 46398 7698
rect 46450 7646 46452 7698
rect 46060 7644 46452 7646
rect 46060 7634 46116 7644
rect 46396 7634 46452 7644
rect 46508 7644 46900 7700
rect 45836 7586 46004 7588
rect 45836 7534 45838 7586
rect 45890 7534 46004 7586
rect 45836 7532 46004 7534
rect 45388 7310 45390 7362
rect 45442 7310 45444 7362
rect 45388 7298 45444 7310
rect 45724 7474 45780 7486
rect 45724 7422 45726 7474
rect 45778 7422 45780 7474
rect 44268 6862 44270 6914
rect 44322 6862 44324 6914
rect 44268 6850 44324 6862
rect 44716 7196 44996 7252
rect 43708 6738 43764 6748
rect 44268 6692 44324 6702
rect 44324 6636 44548 6692
rect 44268 6598 44324 6636
rect 43596 6402 43652 6412
rect 44132 6300 44396 6310
rect 44188 6244 44236 6300
rect 44292 6244 44340 6300
rect 44132 6234 44396 6244
rect 43372 5182 43374 5234
rect 43426 5182 43428 5234
rect 43372 4900 43428 5182
rect 43596 5122 43652 5134
rect 43596 5070 43598 5122
rect 43650 5070 43652 5122
rect 43596 5012 43652 5070
rect 43820 5124 43876 5134
rect 43820 5030 43876 5068
rect 43596 4956 43764 5012
rect 43372 4844 43652 4900
rect 42588 4338 42756 4340
rect 42588 4286 42590 4338
rect 42642 4286 42756 4338
rect 42588 4284 42756 4286
rect 43596 4340 43652 4844
rect 43708 4676 43764 4956
rect 44132 4732 44396 4742
rect 44188 4676 44236 4732
rect 44292 4676 44340 4732
rect 43764 4620 43988 4676
rect 44132 4666 44396 4676
rect 43708 4610 43764 4620
rect 43932 4452 43988 4620
rect 44492 4562 44548 6636
rect 44492 4510 44494 4562
rect 44546 4510 44548 4562
rect 44492 4498 44548 4510
rect 43820 4340 43876 4350
rect 43596 4338 43876 4340
rect 43596 4286 43822 4338
rect 43874 4286 43876 4338
rect 43596 4284 43876 4286
rect 42588 4274 42644 4284
rect 43820 4274 43876 4284
rect 43932 3666 43988 4396
rect 44156 4340 44212 4350
rect 44156 4246 44212 4284
rect 43932 3614 43934 3666
rect 43986 3614 43988 3666
rect 43932 3602 43988 3614
rect 44716 3666 44772 7196
rect 44828 6916 44884 6926
rect 44828 6690 44884 6860
rect 44828 6638 44830 6690
rect 44882 6638 44884 6690
rect 44828 6626 44884 6638
rect 45388 6804 45444 6814
rect 44716 3614 44718 3666
rect 44770 3614 44772 3666
rect 44716 3602 44772 3614
rect 44828 5908 44884 5918
rect 44828 5124 44884 5852
rect 45388 5796 45444 6748
rect 45724 6580 45780 7422
rect 45724 6514 45780 6524
rect 45388 5730 45444 5740
rect 45836 6468 45892 7532
rect 46284 7476 46340 7486
rect 46284 7382 46340 7420
rect 46060 6692 46116 6702
rect 46060 6598 46116 6636
rect 46508 6580 46564 7644
rect 46956 7586 47012 7598
rect 46956 7534 46958 7586
rect 47010 7534 47012 7586
rect 46620 7476 46676 7486
rect 46844 7476 46900 7486
rect 46620 7474 46900 7476
rect 46620 7422 46622 7474
rect 46674 7422 46846 7474
rect 46898 7422 46900 7474
rect 46620 7420 46900 7422
rect 46620 7410 46676 7420
rect 46844 7410 46900 7420
rect 46844 6916 46900 6926
rect 46956 6916 47012 7534
rect 46844 6914 47012 6916
rect 46844 6862 46846 6914
rect 46898 6862 47012 6914
rect 46844 6860 47012 6862
rect 46508 6514 46564 6524
rect 46732 6690 46788 6702
rect 46732 6638 46734 6690
rect 46786 6638 46788 6690
rect 45836 5236 45892 6412
rect 46732 6468 46788 6638
rect 46844 6692 46900 6860
rect 46844 6626 46900 6636
rect 46732 6402 46788 6412
rect 47068 6132 47124 8988
rect 47628 8978 47684 8988
rect 47516 8820 47572 8830
rect 47516 8726 47572 8764
rect 47740 8484 47796 8988
rect 47852 8820 47908 8830
rect 47964 8820 48020 9324
rect 48300 9268 48356 9996
rect 48412 9826 48468 9838
rect 48412 9774 48414 9826
rect 48466 9774 48468 9826
rect 48412 9604 48468 9774
rect 48412 9538 48468 9548
rect 48524 9826 48580 9838
rect 48524 9774 48526 9826
rect 48578 9774 48580 9826
rect 48076 9212 48356 9268
rect 48076 9042 48132 9212
rect 48076 8990 48078 9042
rect 48130 8990 48132 9042
rect 48076 8978 48132 8990
rect 48188 9044 48244 9054
rect 48188 8950 48244 8988
rect 47852 8818 48020 8820
rect 47852 8766 47854 8818
rect 47906 8766 48020 8818
rect 47852 8764 48020 8766
rect 47852 8754 47908 8764
rect 47852 8484 47908 8494
rect 47740 8482 47908 8484
rect 47740 8430 47854 8482
rect 47906 8430 47908 8482
rect 47740 8428 47908 8430
rect 47852 8418 47908 8428
rect 47628 8260 47684 8270
rect 47180 8258 47684 8260
rect 47180 8206 47630 8258
rect 47682 8206 47684 8258
rect 47180 8204 47684 8206
rect 47964 8260 48020 8764
rect 48300 8482 48356 9212
rect 48300 8430 48302 8482
rect 48354 8430 48356 8482
rect 48300 8418 48356 8430
rect 48076 8260 48132 8270
rect 47964 8258 48132 8260
rect 47964 8206 48078 8258
rect 48130 8206 48132 8258
rect 47964 8204 48132 8206
rect 47180 7698 47236 8204
rect 47628 8194 47684 8204
rect 48076 8036 48132 8204
rect 48412 8260 48468 8270
rect 48412 8166 48468 8204
rect 48076 7970 48132 7980
rect 47180 7646 47182 7698
rect 47234 7646 47236 7698
rect 47180 7634 47236 7646
rect 48076 7364 48132 7374
rect 47964 7362 48132 7364
rect 47964 7310 48078 7362
rect 48130 7310 48132 7362
rect 47964 7308 48132 7310
rect 47180 6690 47236 6702
rect 47180 6638 47182 6690
rect 47234 6638 47236 6690
rect 47180 6580 47236 6638
rect 47180 6514 47236 6524
rect 45836 5170 45892 5180
rect 46732 6076 47124 6132
rect 47740 6356 47796 6366
rect 45276 5124 45332 5134
rect 44828 5122 45332 5124
rect 44828 5070 45278 5122
rect 45330 5070 45332 5122
rect 44828 5068 45332 5070
rect 44828 3554 44884 5068
rect 45276 5058 45332 5068
rect 45612 5124 45668 5134
rect 45612 5030 45668 5068
rect 46732 5122 46788 6076
rect 46732 5070 46734 5122
rect 46786 5070 46788 5122
rect 44940 4898 44996 4910
rect 44940 4846 44942 4898
rect 44994 4846 44996 4898
rect 44940 4788 44996 4846
rect 44940 4722 44996 4732
rect 46732 4788 46788 5070
rect 46844 5906 46900 5918
rect 46844 5854 46846 5906
rect 46898 5854 46900 5906
rect 46844 5124 46900 5854
rect 47068 5906 47124 5918
rect 47068 5854 47070 5906
rect 47122 5854 47124 5906
rect 47068 5346 47124 5854
rect 47068 5294 47070 5346
rect 47122 5294 47124 5346
rect 47068 5282 47124 5294
rect 47628 5906 47684 5918
rect 47628 5854 47630 5906
rect 47682 5854 47684 5906
rect 46844 5058 46900 5068
rect 45164 4452 45220 4462
rect 45164 4358 45220 4396
rect 46732 4452 46788 4732
rect 47404 4452 47460 4462
rect 46788 4396 46900 4452
rect 46732 4386 46788 4396
rect 46844 3666 46900 4396
rect 47404 4358 47460 4396
rect 46844 3614 46846 3666
rect 46898 3614 46900 3666
rect 46844 3602 46900 3614
rect 47628 3666 47684 5854
rect 47740 4450 47796 6300
rect 47964 5348 48020 7308
rect 48076 7298 48132 7308
rect 48300 6692 48356 6702
rect 48076 6020 48132 6030
rect 48076 5926 48132 5964
rect 48076 5348 48132 5358
rect 47964 5292 48076 5348
rect 48076 5282 48132 5292
rect 48300 5124 48356 6636
rect 48524 6690 48580 9774
rect 48748 9154 48804 9996
rect 48972 9380 49028 12124
rect 49420 12086 49476 12124
rect 49308 12068 49364 12078
rect 49196 12066 49364 12068
rect 49196 12014 49310 12066
rect 49362 12014 49364 12066
rect 49196 12012 49364 12014
rect 49084 11956 49140 11966
rect 49084 11862 49140 11900
rect 49084 11732 49140 11742
rect 49084 11506 49140 11676
rect 49084 11454 49086 11506
rect 49138 11454 49140 11506
rect 49084 11442 49140 11454
rect 49084 9828 49140 9838
rect 49196 9828 49252 12012
rect 49308 12002 49364 12012
rect 49532 11396 49588 12572
rect 49644 12404 49700 12414
rect 49980 12404 50036 13134
rect 49644 12290 49700 12348
rect 49644 12238 49646 12290
rect 49698 12238 49700 12290
rect 49644 12226 49700 12238
rect 49868 12348 50036 12404
rect 50092 13132 50204 13188
rect 50260 13132 50372 13188
rect 50092 12404 50148 13132
rect 50204 13122 50260 13132
rect 50316 13074 50372 13132
rect 50316 13022 50318 13074
rect 50370 13022 50372 13074
rect 50316 13010 50372 13022
rect 49868 11732 49924 12348
rect 50092 12310 50148 12348
rect 49868 11666 49924 11676
rect 49980 12180 50036 12190
rect 49532 11340 49700 11396
rect 49532 11172 49588 11182
rect 49420 11170 49588 11172
rect 49420 11118 49534 11170
rect 49586 11118 49588 11170
rect 49420 11116 49588 11118
rect 49308 10612 49364 10622
rect 49420 10612 49476 11116
rect 49532 11106 49588 11116
rect 49644 11060 49700 11340
rect 49700 11004 49812 11060
rect 49644 10994 49700 11004
rect 49756 10722 49812 11004
rect 49756 10670 49758 10722
rect 49810 10670 49812 10722
rect 49756 10658 49812 10670
rect 49980 10722 50036 12124
rect 50316 11508 50372 11518
rect 50316 11414 50372 11452
rect 49980 10670 49982 10722
rect 50034 10670 50036 10722
rect 49980 10658 50036 10670
rect 50428 10724 50484 14476
rect 50540 14308 50596 14318
rect 50876 14308 50932 14478
rect 50596 14252 50932 14308
rect 50988 14530 51268 14532
rect 50988 14478 51214 14530
rect 51266 14478 51268 14530
rect 50988 14476 51268 14478
rect 50540 14214 50596 14252
rect 50988 12964 51044 14476
rect 51212 14466 51268 14476
rect 51436 14530 51492 14542
rect 51436 14478 51438 14530
rect 51490 14478 51492 14530
rect 51100 14306 51156 14318
rect 51100 14254 51102 14306
rect 51154 14254 51156 14306
rect 51100 13860 51156 14254
rect 51100 13794 51156 13804
rect 51212 13972 51268 13982
rect 51436 13972 51492 14478
rect 51212 13970 51492 13972
rect 51212 13918 51214 13970
rect 51266 13918 51492 13970
rect 51212 13916 51492 13918
rect 51212 13524 51268 13916
rect 50652 12908 50988 12964
rect 50652 11506 50708 12908
rect 50988 12898 51044 12908
rect 51100 13468 51212 13524
rect 51100 12962 51156 13468
rect 51212 13458 51268 13468
rect 51660 13858 51716 13870
rect 51660 13806 51662 13858
rect 51714 13806 51716 13858
rect 51286 13356 51550 13366
rect 51342 13300 51390 13356
rect 51446 13300 51494 13356
rect 51286 13290 51550 13300
rect 51660 13188 51716 13806
rect 51660 13122 51716 13132
rect 51436 13076 51492 13086
rect 51436 12982 51492 13020
rect 51100 12910 51102 12962
rect 51154 12910 51156 12962
rect 50764 12738 50820 12750
rect 50764 12686 50766 12738
rect 50818 12686 50820 12738
rect 50764 12402 50820 12686
rect 50764 12350 50766 12402
rect 50818 12350 50820 12402
rect 50764 11620 50820 12350
rect 51100 12180 51156 12910
rect 51324 12964 51380 12974
rect 51324 12290 51380 12908
rect 51548 12852 51604 12862
rect 51548 12758 51604 12796
rect 51324 12238 51326 12290
rect 51378 12238 51380 12290
rect 51324 12226 51380 12238
rect 51660 12292 51716 12302
rect 51660 12198 51716 12236
rect 51100 12086 51156 12124
rect 51548 12068 51604 12078
rect 51548 11974 51604 12012
rect 51286 11788 51550 11798
rect 51342 11732 51390 11788
rect 51446 11732 51494 11788
rect 51286 11722 51550 11732
rect 50764 11554 50820 11564
rect 50652 11454 50654 11506
rect 50706 11454 50708 11506
rect 50652 11060 50708 11454
rect 51772 11508 51828 15092
rect 53452 14868 53508 14878
rect 51772 11414 51828 11452
rect 51884 14756 51940 14766
rect 50428 10668 50596 10724
rect 49308 10610 49476 10612
rect 49308 10558 49310 10610
rect 49362 10558 49476 10610
rect 49308 10556 49476 10558
rect 49644 10612 49700 10622
rect 49308 10276 49364 10556
rect 49308 10210 49364 10220
rect 49532 10498 49588 10510
rect 49532 10446 49534 10498
rect 49586 10446 49588 10498
rect 49532 10052 49588 10446
rect 49084 9826 49252 9828
rect 49084 9774 49086 9826
rect 49138 9774 49252 9826
rect 49084 9772 49252 9774
rect 49308 9996 49588 10052
rect 49644 10050 49700 10556
rect 50428 10500 50484 10510
rect 50428 10406 50484 10444
rect 49644 9998 49646 10050
rect 49698 9998 49700 10050
rect 49308 9826 49364 9996
rect 49644 9986 49700 9998
rect 49980 10052 50036 10062
rect 49980 9938 50036 9996
rect 49980 9886 49982 9938
rect 50034 9886 50036 9938
rect 49308 9774 49310 9826
rect 49362 9774 49364 9826
rect 49084 9762 49140 9772
rect 49308 9762 49364 9774
rect 49532 9828 49588 9838
rect 49532 9714 49588 9772
rect 49532 9662 49534 9714
rect 49586 9662 49588 9714
rect 49532 9650 49588 9662
rect 49868 9716 49924 9726
rect 48748 9102 48750 9154
rect 48802 9102 48804 9154
rect 48748 9090 48804 9102
rect 48860 9324 49028 9380
rect 48748 8932 48804 8942
rect 48748 8484 48804 8876
rect 48860 8596 48916 9324
rect 48972 9154 49028 9166
rect 48972 9102 48974 9154
rect 49026 9102 49028 9154
rect 48972 9044 49028 9102
rect 48972 8978 49028 8988
rect 49084 8820 49140 8830
rect 49084 8818 49364 8820
rect 49084 8766 49086 8818
rect 49138 8766 49364 8818
rect 49084 8764 49364 8766
rect 49084 8754 49140 8764
rect 48860 8540 49140 8596
rect 48748 8428 48916 8484
rect 48748 8260 48804 8270
rect 48748 8166 48804 8204
rect 48860 7698 48916 8428
rect 49084 8370 49140 8540
rect 49084 8318 49086 8370
rect 49138 8318 49140 8370
rect 49084 8306 49140 8318
rect 48860 7646 48862 7698
rect 48914 7646 48916 7698
rect 48524 6638 48526 6690
rect 48578 6638 48580 6690
rect 48524 6626 48580 6638
rect 48748 6690 48804 6702
rect 48748 6638 48750 6690
rect 48802 6638 48804 6690
rect 48748 6356 48804 6638
rect 48860 6580 48916 7646
rect 48972 8034 49028 8046
rect 48972 7982 48974 8034
rect 49026 7982 49028 8034
rect 48972 6916 49028 7982
rect 48972 6860 49252 6916
rect 48972 6692 49028 6702
rect 48972 6598 49028 6636
rect 48860 6514 48916 6524
rect 48748 5236 48804 6300
rect 48860 5906 48916 5918
rect 48860 5854 48862 5906
rect 48914 5854 48916 5906
rect 48860 5348 48916 5854
rect 48972 5908 49028 5918
rect 48972 5814 49028 5852
rect 49084 5906 49140 5918
rect 49084 5854 49086 5906
rect 49138 5854 49140 5906
rect 48860 5282 48916 5292
rect 49084 5460 49140 5854
rect 49196 5906 49252 6860
rect 49196 5854 49198 5906
rect 49250 5854 49252 5906
rect 49196 5842 49252 5854
rect 47964 5122 48356 5124
rect 47964 5070 48302 5122
rect 48354 5070 48356 5122
rect 47964 5068 48356 5070
rect 47964 4562 48020 5068
rect 47964 4510 47966 4562
rect 48018 4510 48020 4562
rect 47964 4498 48020 4510
rect 47740 4398 47742 4450
rect 47794 4398 47796 4450
rect 47740 4386 47796 4398
rect 48076 4228 48132 4238
rect 48076 4134 48132 4172
rect 47628 3614 47630 3666
rect 47682 3614 47684 3666
rect 47628 3602 47684 3614
rect 48188 3666 48244 5068
rect 48300 5058 48356 5068
rect 48524 5234 48804 5236
rect 48524 5182 48750 5234
rect 48802 5182 48804 5234
rect 48524 5180 48804 5182
rect 48188 3614 48190 3666
rect 48242 3614 48244 3666
rect 48188 3602 48244 3614
rect 44828 3502 44830 3554
rect 44882 3502 44884 3554
rect 44828 3490 44884 3502
rect 48524 3554 48580 5180
rect 48748 5170 48804 5180
rect 48972 4900 49028 4910
rect 49084 4900 49140 5404
rect 49196 5348 49252 5358
rect 49196 5254 49252 5292
rect 49308 5236 49364 8764
rect 49532 6580 49588 6590
rect 49532 5906 49588 6524
rect 49868 6244 49924 9660
rect 49980 8932 50036 9886
rect 50428 9268 50484 9278
rect 50540 9268 50596 10668
rect 50652 10500 50708 11004
rect 50652 10434 50708 10444
rect 51660 11394 51716 11406
rect 51660 11342 51662 11394
rect 51714 11342 51716 11394
rect 51286 10220 51550 10230
rect 51342 10164 51390 10220
rect 51446 10164 51494 10220
rect 51286 10154 51550 10164
rect 51660 9940 51716 11342
rect 51660 9874 51716 9884
rect 51772 10722 51828 10734
rect 51772 10670 51774 10722
rect 51826 10670 51828 10722
rect 50428 9266 51044 9268
rect 50428 9214 50430 9266
rect 50482 9214 51044 9266
rect 50428 9212 51044 9214
rect 50428 9202 50484 9212
rect 49980 8866 50036 8876
rect 50316 8372 50372 8382
rect 50652 8372 50708 9212
rect 50316 8370 50708 8372
rect 50316 8318 50318 8370
rect 50370 8318 50654 8370
rect 50706 8318 50708 8370
rect 50316 8316 50708 8318
rect 50316 8306 50372 8316
rect 50652 8306 50708 8316
rect 50764 9044 50820 9054
rect 50764 8260 50820 8988
rect 50988 9042 51044 9212
rect 50988 8990 50990 9042
rect 51042 8990 51044 9042
rect 50988 8978 51044 8990
rect 51324 8932 51380 8942
rect 51324 8838 51380 8876
rect 51772 8932 51828 10670
rect 51772 8866 51828 8876
rect 51286 8652 51550 8662
rect 51342 8596 51390 8652
rect 51446 8596 51494 8652
rect 51286 8586 51550 8596
rect 50876 8260 50932 8270
rect 50764 8258 50932 8260
rect 50764 8206 50878 8258
rect 50930 8206 50932 8258
rect 50764 8204 50932 8206
rect 50876 8194 50932 8204
rect 51548 8148 51604 8158
rect 51548 8146 51716 8148
rect 51548 8094 51550 8146
rect 51602 8094 51716 8146
rect 51548 8092 51716 8094
rect 51548 8082 51604 8092
rect 51286 7084 51550 7094
rect 51342 7028 51390 7084
rect 51446 7028 51494 7084
rect 51286 7018 51550 7028
rect 51100 6802 51156 6814
rect 51100 6750 51102 6802
rect 51154 6750 51156 6802
rect 50764 6690 50820 6702
rect 50764 6638 50766 6690
rect 50818 6638 50820 6690
rect 50092 6468 50148 6478
rect 50092 6466 50372 6468
rect 50092 6414 50094 6466
rect 50146 6414 50372 6466
rect 50092 6412 50372 6414
rect 50092 6402 50148 6412
rect 50316 6244 50372 6412
rect 49868 6188 50148 6244
rect 50092 6020 50148 6188
rect 50092 5926 50148 5964
rect 49532 5854 49534 5906
rect 49586 5854 49588 5906
rect 49532 5348 49588 5854
rect 50316 5906 50372 6188
rect 50652 6132 50708 6142
rect 50764 6132 50820 6638
rect 51100 6692 51156 6750
rect 51100 6626 51156 6636
rect 51548 6692 51604 6702
rect 51660 6692 51716 8092
rect 51604 6636 51716 6692
rect 51548 6626 51604 6636
rect 51324 6580 51380 6590
rect 50652 6130 50764 6132
rect 50652 6078 50654 6130
rect 50706 6078 50764 6130
rect 50652 6076 50764 6078
rect 50652 6066 50708 6076
rect 50764 6038 50820 6076
rect 50988 6244 51044 6254
rect 50988 6018 51044 6188
rect 51324 6130 51380 6524
rect 51884 6244 51940 14700
rect 53452 14642 53508 14812
rect 53452 14590 53454 14642
rect 53506 14590 53508 14642
rect 53452 14578 53508 14590
rect 53004 14530 53060 14542
rect 53004 14478 53006 14530
rect 53058 14478 53060 14530
rect 52108 14308 52164 14318
rect 52108 14214 52164 14252
rect 52556 14308 52612 14318
rect 53004 14308 53060 14478
rect 52556 14306 52836 14308
rect 52556 14254 52558 14306
rect 52610 14254 52836 14306
rect 52556 14252 52836 14254
rect 52556 14242 52612 14252
rect 52556 13746 52612 13758
rect 52556 13694 52558 13746
rect 52610 13694 52612 13746
rect 52556 12964 52612 13694
rect 51996 12852 52052 12862
rect 51996 12758 52052 12796
rect 52556 12402 52612 12908
rect 52668 13188 52724 13198
rect 52668 12964 52724 13132
rect 52780 13076 52836 14252
rect 53004 14242 53060 14252
rect 53228 14530 53284 14542
rect 53228 14478 53230 14530
rect 53282 14478 53284 14530
rect 53228 14084 53284 14478
rect 53228 14018 53284 14028
rect 52892 13636 52948 13646
rect 52892 13634 53060 13636
rect 52892 13582 52894 13634
rect 52946 13582 53060 13634
rect 52892 13580 53060 13582
rect 52892 13570 52948 13580
rect 52892 13076 52948 13086
rect 52780 13074 52948 13076
rect 52780 13022 52894 13074
rect 52946 13022 52948 13074
rect 52780 13020 52948 13022
rect 52892 13010 52948 13020
rect 53004 12964 53060 13580
rect 53116 13524 53172 13534
rect 53116 13186 53172 13468
rect 53116 13134 53118 13186
rect 53170 13134 53172 13186
rect 53116 13122 53172 13134
rect 53564 13076 53620 17052
rect 53676 16212 53732 16222
rect 53676 16098 53732 16156
rect 53676 16046 53678 16098
rect 53730 16046 53732 16098
rect 53676 16034 53732 16046
rect 53676 15316 53732 15326
rect 53788 15316 53844 18060
rect 54012 17892 54068 17902
rect 53900 16996 53956 17034
rect 53900 16930 53956 16940
rect 53676 15314 53844 15316
rect 53676 15262 53678 15314
rect 53730 15262 53844 15314
rect 53676 15260 53844 15262
rect 53676 15250 53732 15260
rect 53788 15204 53844 15260
rect 53788 15138 53844 15148
rect 53900 16772 53956 16782
rect 53900 15202 53956 16716
rect 54012 16322 54068 17836
rect 54236 17666 54292 18284
rect 54236 17614 54238 17666
rect 54290 17614 54292 17666
rect 54236 17444 54292 17614
rect 54236 17378 54292 17388
rect 54460 16660 54516 18284
rect 54572 17892 54628 17902
rect 54572 17666 54628 17836
rect 55020 17668 55076 18732
rect 54572 17614 54574 17666
rect 54626 17614 54628 17666
rect 54572 17602 54628 17614
rect 54908 17612 55076 17668
rect 55132 18564 55188 18574
rect 54796 17332 54852 17342
rect 54451 16604 54516 16660
rect 54684 17276 54796 17332
rect 54451 16548 54507 16604
rect 54451 16492 54516 16548
rect 54012 16270 54014 16322
rect 54066 16270 54068 16322
rect 54012 16258 54068 16270
rect 54348 16100 54404 16110
rect 54124 15316 54180 15326
rect 54348 15316 54404 16044
rect 54124 15314 54404 15316
rect 54124 15262 54126 15314
rect 54178 15262 54404 15314
rect 54124 15260 54404 15262
rect 54124 15250 54180 15260
rect 53900 15150 53902 15202
rect 53954 15150 53956 15202
rect 53900 15138 53956 15150
rect 54012 15204 54068 15214
rect 53900 14980 53956 14990
rect 53564 13010 53620 13020
rect 53788 14308 53844 14318
rect 53788 13076 53844 14252
rect 53676 12964 53732 12974
rect 52668 12962 52836 12964
rect 52668 12910 52670 12962
rect 52722 12910 52836 12962
rect 52668 12908 52836 12910
rect 53004 12908 53172 12964
rect 52668 12898 52724 12908
rect 52780 12852 52836 12908
rect 52780 12796 53060 12852
rect 52556 12350 52558 12402
rect 52610 12350 52612 12402
rect 52556 12338 52612 12350
rect 53004 12402 53060 12796
rect 53004 12350 53006 12402
rect 53058 12350 53060 12402
rect 53004 12338 53060 12350
rect 52108 12292 52164 12302
rect 52108 12198 52164 12236
rect 53116 11620 53172 12908
rect 53676 12870 53732 12908
rect 53228 12852 53284 12862
rect 53228 12738 53284 12796
rect 53228 12686 53230 12738
rect 53282 12686 53284 12738
rect 53228 12674 53284 12686
rect 53340 12850 53396 12862
rect 53340 12798 53342 12850
rect 53394 12798 53396 12850
rect 53340 12740 53396 12798
rect 53116 11554 53172 11564
rect 53228 11732 53284 11742
rect 53228 11396 53284 11676
rect 52108 11284 52164 11294
rect 51996 11282 52164 11284
rect 51996 11230 52110 11282
rect 52162 11230 52164 11282
rect 51996 11228 52164 11230
rect 51996 10610 52052 11228
rect 52108 11218 52164 11228
rect 51996 10558 51998 10610
rect 52050 10558 52052 10610
rect 51996 10546 52052 10558
rect 52892 10610 52948 10622
rect 52892 10558 52894 10610
rect 52946 10558 52948 10610
rect 52892 9042 52948 10558
rect 53228 9044 53284 11340
rect 52892 8990 52894 9042
rect 52946 8990 52948 9042
rect 52108 8930 52164 8942
rect 52108 8878 52110 8930
rect 52162 8878 52164 8930
rect 52108 8372 52164 8878
rect 52108 8306 52164 8316
rect 52892 8260 52948 8990
rect 52892 8194 52948 8204
rect 53004 9042 53284 9044
rect 53004 8990 53230 9042
rect 53282 8990 53284 9042
rect 53004 8988 53284 8990
rect 53004 8372 53060 8988
rect 53228 8978 53284 8988
rect 52892 8036 52948 8046
rect 53004 8036 53060 8316
rect 52892 8034 53060 8036
rect 52892 7982 52894 8034
rect 52946 7982 53060 8034
rect 52892 7980 53060 7982
rect 52892 7970 52948 7980
rect 52780 6916 52836 6926
rect 52780 6822 52836 6860
rect 53228 6804 53284 6814
rect 53340 6804 53396 12684
rect 53788 12066 53844 13020
rect 53788 12014 53790 12066
rect 53842 12014 53844 12066
rect 53788 11956 53844 12014
rect 53788 11890 53844 11900
rect 53900 11732 53956 14924
rect 54012 13748 54068 15148
rect 54460 14756 54516 16492
rect 54684 16436 54740 17276
rect 54796 17266 54852 17276
rect 54684 16380 54852 16436
rect 54572 16324 54628 16334
rect 54572 16210 54628 16268
rect 54572 16158 54574 16210
rect 54626 16158 54628 16210
rect 54572 14980 54628 16158
rect 54684 16212 54740 16222
rect 54684 15426 54740 16156
rect 54796 15540 54852 16380
rect 54908 16100 54964 17612
rect 55132 17554 55188 18508
rect 55132 17502 55134 17554
rect 55186 17502 55188 17554
rect 55132 17490 55188 17502
rect 55020 17442 55076 17454
rect 55020 17390 55022 17442
rect 55074 17390 55076 17442
rect 55020 16436 55076 17390
rect 55020 16370 55076 16380
rect 55244 17444 55300 17454
rect 55244 16100 55300 17388
rect 55356 17332 55412 17342
rect 55412 17276 55524 17332
rect 55356 17266 55412 17276
rect 55468 17106 55524 17276
rect 55468 17054 55470 17106
rect 55522 17054 55524 17106
rect 55468 17042 55524 17054
rect 55580 16772 55636 21308
rect 55692 21298 55748 21308
rect 55692 20802 55748 20814
rect 55692 20750 55694 20802
rect 55746 20750 55748 20802
rect 55692 20692 55748 20750
rect 55692 20626 55748 20636
rect 55804 20244 55860 21532
rect 56028 21476 56084 21646
rect 56028 21410 56084 21420
rect 56476 22146 56532 22158
rect 56476 22094 56478 22146
rect 56530 22094 56532 22146
rect 56476 20916 56532 22094
rect 56700 21476 56756 21486
rect 56700 21382 56756 21420
rect 56028 20914 56532 20916
rect 56028 20862 56478 20914
rect 56530 20862 56532 20914
rect 56028 20860 56532 20862
rect 55916 20244 55972 20254
rect 55804 20242 55972 20244
rect 55804 20190 55918 20242
rect 55970 20190 55972 20242
rect 55804 20188 55972 20190
rect 55916 20178 55972 20188
rect 56028 19348 56084 20860
rect 56476 20850 56532 20860
rect 55692 19292 56084 19348
rect 56140 20692 56196 20702
rect 55692 18564 55748 19292
rect 55692 18508 55972 18564
rect 55692 17666 55748 18508
rect 55692 17614 55694 17666
rect 55746 17614 55748 17666
rect 55692 17602 55748 17614
rect 55804 18338 55860 18350
rect 55804 18286 55806 18338
rect 55858 18286 55860 18338
rect 55580 16706 55636 16716
rect 55692 16882 55748 16894
rect 55692 16830 55694 16882
rect 55746 16830 55748 16882
rect 54908 16006 54964 16044
rect 55132 16044 55300 16100
rect 55356 16658 55412 16670
rect 55356 16606 55358 16658
rect 55410 16606 55412 16658
rect 55356 16100 55412 16606
rect 55020 15988 55076 15998
rect 55020 15894 55076 15932
rect 54796 15474 54852 15484
rect 54684 15374 54686 15426
rect 54738 15374 54740 15426
rect 54684 15362 54740 15374
rect 55132 15316 55188 16044
rect 55356 16034 55412 16044
rect 55468 16436 55524 16446
rect 55244 15876 55300 15886
rect 55244 15874 55412 15876
rect 55244 15822 55246 15874
rect 55298 15822 55412 15874
rect 55244 15820 55412 15822
rect 55244 15810 55300 15820
rect 55244 15540 55300 15550
rect 55244 15446 55300 15484
rect 55132 15148 55188 15260
rect 54572 14914 54628 14924
rect 54796 15092 55188 15148
rect 54460 14700 54740 14756
rect 54460 14530 54516 14542
rect 54460 14478 54462 14530
rect 54514 14478 54516 14530
rect 54348 13748 54404 13758
rect 54012 13746 54404 13748
rect 54012 13694 54350 13746
rect 54402 13694 54404 13746
rect 54012 13692 54404 13694
rect 54348 13682 54404 13692
rect 54460 13524 54516 14478
rect 54572 14308 54628 14318
rect 54572 14214 54628 14252
rect 54684 13748 54740 14700
rect 54684 13682 54740 13692
rect 54796 13746 54852 15092
rect 55132 14868 55188 14878
rect 55020 14812 55132 14868
rect 55020 14418 55076 14812
rect 55132 14802 55188 14812
rect 55020 14366 55022 14418
rect 55074 14366 55076 14418
rect 55020 14354 55076 14366
rect 55356 14420 55412 15820
rect 55468 15148 55524 16380
rect 55692 16324 55748 16830
rect 55692 16258 55748 16268
rect 55580 16212 55636 16222
rect 55580 16118 55636 16156
rect 55804 16098 55860 18286
rect 55916 16994 55972 18508
rect 56140 17554 56196 20636
rect 56812 20692 56868 23660
rect 56924 23268 56980 23884
rect 56924 23154 56980 23212
rect 56924 23102 56926 23154
rect 56978 23102 56980 23154
rect 56924 23090 56980 23102
rect 57036 23380 57092 24444
rect 57148 24498 57204 24510
rect 57148 24446 57150 24498
rect 57202 24446 57204 24498
rect 57148 23380 57204 24446
rect 57708 23940 57764 23950
rect 57596 23716 57652 23726
rect 57596 23622 57652 23660
rect 57148 23324 57428 23380
rect 57036 23042 57092 23324
rect 57036 22990 57038 23042
rect 57090 22990 57092 23042
rect 57036 22978 57092 22990
rect 57260 22930 57316 22942
rect 57260 22878 57262 22930
rect 57314 22878 57316 22930
rect 57260 21588 57316 22878
rect 57372 22260 57428 23324
rect 57484 22260 57540 22270
rect 57372 22258 57540 22260
rect 57372 22206 57486 22258
rect 57538 22206 57540 22258
rect 57372 22204 57540 22206
rect 57484 22194 57540 22204
rect 57708 21812 57764 23884
rect 57932 23938 57988 23950
rect 57932 23886 57934 23938
rect 57986 23886 57988 23938
rect 57932 23604 57988 23886
rect 57932 23538 57988 23548
rect 58439 23548 58703 23558
rect 58495 23492 58543 23548
rect 58599 23492 58647 23548
rect 58439 23482 58703 23492
rect 58439 21980 58703 21990
rect 58495 21924 58543 21980
rect 58599 21924 58647 21980
rect 58439 21914 58703 21924
rect 57708 21756 58212 21812
rect 57708 21698 57764 21756
rect 57708 21646 57710 21698
rect 57762 21646 57764 21698
rect 57708 21634 57764 21646
rect 57932 21588 57988 21598
rect 57260 21586 57428 21588
rect 57260 21534 57262 21586
rect 57314 21534 57428 21586
rect 57260 21532 57428 21534
rect 57260 21522 57316 21532
rect 57372 21252 57428 21532
rect 57372 21196 57764 21252
rect 57708 20802 57764 21196
rect 57708 20750 57710 20802
rect 57762 20750 57764 20802
rect 57708 20738 57764 20750
rect 57932 20802 57988 21532
rect 57932 20750 57934 20802
rect 57986 20750 57988 20802
rect 57932 20738 57988 20750
rect 58044 21474 58100 21486
rect 58044 21422 58046 21474
rect 58098 21422 58100 21474
rect 56812 20690 57092 20692
rect 56812 20638 56814 20690
rect 56866 20638 57092 20690
rect 56812 20636 57092 20638
rect 56812 20626 56868 20636
rect 57036 20132 57092 20636
rect 57372 20580 57428 20590
rect 57372 20578 57540 20580
rect 57372 20526 57374 20578
rect 57426 20526 57540 20578
rect 57372 20524 57540 20526
rect 57372 20514 57428 20524
rect 57036 20076 57428 20132
rect 56924 20020 56980 20030
rect 56364 20018 56980 20020
rect 56364 19966 56926 20018
rect 56978 19966 56980 20018
rect 56364 19964 56980 19966
rect 56140 17502 56142 17554
rect 56194 17502 56196 17554
rect 56140 17490 56196 17502
rect 56252 19122 56308 19134
rect 56252 19070 56254 19122
rect 56306 19070 56308 19122
rect 55916 16942 55918 16994
rect 55970 16942 55972 16994
rect 55916 16930 55972 16942
rect 55804 16046 55806 16098
rect 55858 16046 55860 16098
rect 55804 16034 55860 16046
rect 56140 16322 56196 16334
rect 56140 16270 56142 16322
rect 56194 16270 56196 16322
rect 55804 15202 55860 15214
rect 55804 15150 55806 15202
rect 55858 15150 55860 15202
rect 55804 15148 55860 15150
rect 55468 15092 55636 15148
rect 55356 14354 55412 14364
rect 54796 13694 54798 13746
rect 54850 13694 54852 13746
rect 54796 13682 54852 13694
rect 55244 14084 55300 14094
rect 55020 13524 55076 13534
rect 54460 13522 55076 13524
rect 54460 13470 55022 13522
rect 55074 13470 55076 13522
rect 54460 13468 55076 13470
rect 54908 13188 54964 13198
rect 54908 13074 54964 13132
rect 54908 13022 54910 13074
rect 54962 13022 54964 13074
rect 54460 12964 54516 12974
rect 54460 12870 54516 12908
rect 54012 12740 54068 12750
rect 54012 12646 54068 12684
rect 54908 12404 54964 13022
rect 55020 12964 55076 13468
rect 55132 12964 55188 12974
rect 55020 12908 55132 12964
rect 55132 12898 55188 12908
rect 55244 12962 55300 14028
rect 55356 13748 55412 13758
rect 55356 13654 55412 13692
rect 55468 13076 55524 13114
rect 55468 13010 55524 13020
rect 55244 12910 55246 12962
rect 55298 12910 55300 12962
rect 55244 12898 55300 12910
rect 55468 12740 55524 12750
rect 54572 12348 54908 12404
rect 53900 11666 53956 11676
rect 54236 12178 54292 12190
rect 54236 12126 54238 12178
rect 54290 12126 54292 12178
rect 53564 11620 53620 11630
rect 53564 11508 53620 11564
rect 54012 11508 54068 11518
rect 54236 11508 54292 12126
rect 53564 11506 54236 11508
rect 53564 11454 53566 11506
rect 53618 11454 54014 11506
rect 54066 11454 54236 11506
rect 53564 11452 54236 11454
rect 53564 11442 53620 11452
rect 54012 11442 54068 11452
rect 54236 11414 54292 11452
rect 54572 11172 54628 12348
rect 54908 12338 54964 12348
rect 55356 12404 55412 12414
rect 55356 12310 55412 12348
rect 54684 12178 54740 12190
rect 54684 12126 54686 12178
rect 54738 12126 54740 12178
rect 54684 11396 54740 12126
rect 54796 12180 54852 12190
rect 54796 12086 54852 12124
rect 54908 12180 54964 12190
rect 55468 12180 55524 12684
rect 55580 12402 55636 15092
rect 55692 15092 55860 15148
rect 55692 13748 55748 15092
rect 55804 14532 55860 14542
rect 55804 13970 55860 14476
rect 56140 14084 56196 16270
rect 56252 14868 56308 19070
rect 56252 14802 56308 14812
rect 56140 14018 56196 14028
rect 55804 13918 55806 13970
rect 55858 13918 55860 13970
rect 55804 13906 55860 13918
rect 55916 13972 55972 13982
rect 55916 13878 55972 13916
rect 56028 13748 56084 13758
rect 55692 13188 55748 13692
rect 55692 13122 55748 13132
rect 55804 13746 56084 13748
rect 55804 13694 56030 13746
rect 56082 13694 56084 13746
rect 55804 13692 56084 13694
rect 55804 13186 55860 13692
rect 56028 13682 56084 13692
rect 56364 13300 56420 19964
rect 56924 19954 56980 19964
rect 57372 17778 57428 20076
rect 57484 19124 57540 20524
rect 57708 20132 57764 20142
rect 57708 20038 57764 20076
rect 58044 19236 58100 21422
rect 58156 20802 58212 21756
rect 58156 20750 58158 20802
rect 58210 20750 58212 20802
rect 58156 20738 58212 20750
rect 58439 20412 58703 20422
rect 58495 20356 58543 20412
rect 58599 20356 58647 20412
rect 58439 20346 58703 20356
rect 58156 19236 58212 19246
rect 58100 19234 58212 19236
rect 58100 19182 58158 19234
rect 58210 19182 58212 19234
rect 58100 19180 58212 19182
rect 58044 19142 58100 19180
rect 58156 19170 58212 19180
rect 57596 19124 57652 19134
rect 57484 19122 57652 19124
rect 57484 19070 57598 19122
rect 57650 19070 57652 19122
rect 57484 19068 57652 19070
rect 57484 18788 57540 19068
rect 57596 19058 57652 19068
rect 58439 18844 58703 18854
rect 58495 18788 58543 18844
rect 58599 18788 58647 18844
rect 58439 18778 58703 18788
rect 57484 18722 57540 18732
rect 57372 17726 57374 17778
rect 57426 17726 57428 17778
rect 57372 17714 57428 17726
rect 57036 17444 57092 17454
rect 56476 16884 56532 16894
rect 56476 15148 56532 16828
rect 57036 16882 57092 17388
rect 58439 17276 58703 17286
rect 58495 17220 58543 17276
rect 58599 17220 58647 17276
rect 58439 17210 58703 17220
rect 58156 17108 58212 17118
rect 57036 16830 57038 16882
rect 57090 16830 57092 16882
rect 57036 16818 57092 16830
rect 57708 16994 57764 17006
rect 57708 16942 57710 16994
rect 57762 16942 57764 16994
rect 56924 16772 56980 16782
rect 56924 16678 56980 16716
rect 57148 16660 57204 16670
rect 57148 15314 57204 16604
rect 57148 15262 57150 15314
rect 57202 15262 57204 15314
rect 57148 15250 57204 15262
rect 57260 16658 57316 16670
rect 57260 16606 57262 16658
rect 57314 16606 57316 16658
rect 56476 15092 56644 15148
rect 56476 14532 56532 14542
rect 56476 14438 56532 14476
rect 56140 13244 56420 13300
rect 55804 13134 55806 13186
rect 55858 13134 55860 13186
rect 55580 12350 55582 12402
rect 55634 12350 55636 12402
rect 55580 12338 55636 12350
rect 55804 13076 55860 13134
rect 55804 12402 55860 13020
rect 56028 13188 56084 13198
rect 56028 12962 56084 13132
rect 56028 12910 56030 12962
rect 56082 12910 56084 12962
rect 56028 12898 56084 12910
rect 56028 12740 56084 12750
rect 55804 12350 55806 12402
rect 55858 12350 55860 12402
rect 55804 12338 55860 12350
rect 55916 12628 55972 12638
rect 55692 12292 55748 12302
rect 55692 12198 55748 12236
rect 54908 12178 55076 12180
rect 54908 12126 54910 12178
rect 54962 12126 55076 12178
rect 54908 12124 55076 12126
rect 55468 12124 55636 12180
rect 54908 12114 54964 12124
rect 55020 11956 55076 12124
rect 55020 11396 55076 11900
rect 55244 11956 55300 11966
rect 55244 11508 55300 11900
rect 55132 11396 55188 11406
rect 54684 11340 54852 11396
rect 55020 11340 55132 11396
rect 54684 11172 54740 11182
rect 54572 11170 54740 11172
rect 54572 11118 54686 11170
rect 54738 11118 54740 11170
rect 54572 11116 54740 11118
rect 54684 11106 54740 11116
rect 54684 10498 54740 10510
rect 54684 10446 54686 10498
rect 54738 10446 54740 10498
rect 54236 10388 54292 10398
rect 54684 10388 54740 10446
rect 54236 10294 54292 10332
rect 54460 10386 54740 10388
rect 54460 10334 54686 10386
rect 54738 10334 54740 10386
rect 54460 10332 54740 10334
rect 54348 9380 54404 9390
rect 54460 9380 54516 10332
rect 54684 10294 54740 10332
rect 54684 9940 54740 9950
rect 54572 9604 54628 9614
rect 54572 9510 54628 9548
rect 54404 9324 54516 9380
rect 54348 9314 54404 9324
rect 54684 9044 54740 9884
rect 54796 9716 54852 11340
rect 54908 11284 54964 11294
rect 54908 11282 55076 11284
rect 54908 11230 54910 11282
rect 54962 11230 55076 11282
rect 54908 11228 55076 11230
rect 54908 11218 54964 11228
rect 54908 9716 54964 9726
rect 54796 9660 54908 9716
rect 54908 9622 54964 9660
rect 54796 9044 54852 9054
rect 54684 8988 54796 9044
rect 53564 8932 53620 8942
rect 53620 8876 53844 8932
rect 53564 8838 53620 8876
rect 53788 8258 53844 8876
rect 53788 8206 53790 8258
rect 53842 8206 53844 8258
rect 53788 8194 53844 8206
rect 53284 6748 53396 6804
rect 54012 8146 54068 8158
rect 54012 8094 54014 8146
rect 54066 8094 54068 8146
rect 53228 6738 53284 6748
rect 52108 6692 52164 6702
rect 51996 6468 52052 6478
rect 51996 6374 52052 6412
rect 51324 6078 51326 6130
rect 51378 6078 51380 6130
rect 51324 6066 51380 6078
rect 51660 6188 51884 6244
rect 51660 6130 51716 6188
rect 51884 6178 51940 6188
rect 51660 6078 51662 6130
rect 51714 6078 51716 6130
rect 51660 6066 51716 6078
rect 50988 5966 50990 6018
rect 51042 5966 51044 6018
rect 50988 5954 51044 5966
rect 51100 6020 51156 6030
rect 51100 5926 51156 5964
rect 52108 6018 52164 6636
rect 52668 6580 52724 6590
rect 52668 6486 52724 6524
rect 52780 6466 52836 6478
rect 52780 6414 52782 6466
rect 52834 6414 52836 6466
rect 52220 6132 52276 6142
rect 52220 6038 52276 6076
rect 52780 6132 52836 6414
rect 52780 6066 52836 6076
rect 53900 6468 53956 6478
rect 52108 5966 52110 6018
rect 52162 5966 52164 6018
rect 52108 5954 52164 5966
rect 50316 5854 50318 5906
rect 50370 5854 50372 5906
rect 50316 5842 50372 5854
rect 53900 5794 53956 6412
rect 54012 6130 54068 8094
rect 54684 8146 54740 8988
rect 54796 8978 54852 8988
rect 54908 8484 54964 8494
rect 54796 8372 54852 8382
rect 54796 8258 54852 8316
rect 54796 8206 54798 8258
rect 54850 8206 54852 8258
rect 54796 8194 54852 8206
rect 54684 8094 54686 8146
rect 54738 8094 54740 8146
rect 54684 8082 54740 8094
rect 54908 6690 54964 8428
rect 55020 8036 55076 11228
rect 55132 10386 55188 11340
rect 55244 10834 55300 11452
rect 55468 11172 55524 11182
rect 55468 11078 55524 11116
rect 55244 10782 55246 10834
rect 55298 10782 55300 10834
rect 55244 10770 55300 10782
rect 55468 10836 55524 10846
rect 55132 10334 55134 10386
rect 55186 10334 55188 10386
rect 55132 10322 55188 10334
rect 55468 10388 55524 10780
rect 55580 10722 55636 12124
rect 55916 11788 55972 12572
rect 55804 11732 55972 11788
rect 55804 10834 55860 11732
rect 55916 11396 55972 11406
rect 55916 11302 55972 11340
rect 55804 10782 55806 10834
rect 55858 10782 55860 10834
rect 55804 10770 55860 10782
rect 56028 10834 56084 12684
rect 56028 10782 56030 10834
rect 56082 10782 56084 10834
rect 56028 10770 56084 10782
rect 56140 10834 56196 13244
rect 56588 13074 56644 15092
rect 57260 14532 57316 16606
rect 57596 16660 57652 16670
rect 57596 16566 57652 16604
rect 57372 16100 57428 16110
rect 57372 16006 57428 16044
rect 57708 15148 57764 16942
rect 57932 16884 57988 16894
rect 57932 16790 57988 16828
rect 58156 16882 58212 17052
rect 58156 16830 58158 16882
rect 58210 16830 58212 16882
rect 58156 16818 58212 16830
rect 58044 16660 58100 16670
rect 58044 15426 58100 16604
rect 58439 15708 58703 15718
rect 58495 15652 58543 15708
rect 58599 15652 58647 15708
rect 58439 15642 58703 15652
rect 58044 15374 58046 15426
rect 58098 15374 58100 15426
rect 58044 15362 58100 15374
rect 57708 15092 57876 15148
rect 57260 14466 57316 14476
rect 57036 14420 57092 14430
rect 57036 14326 57092 14364
rect 57596 13746 57652 13758
rect 57596 13694 57598 13746
rect 57650 13694 57652 13746
rect 57260 13634 57316 13646
rect 57260 13582 57262 13634
rect 57314 13582 57316 13634
rect 57260 13188 57316 13582
rect 57260 13122 57316 13132
rect 56588 13022 56590 13074
rect 56642 13022 56644 13074
rect 56588 13010 56644 13022
rect 56700 13076 56756 13086
rect 56476 12964 56532 13002
rect 56476 12898 56532 12908
rect 56700 12962 56756 13020
rect 57260 12964 57316 12974
rect 56700 12910 56702 12962
rect 56754 12910 56756 12962
rect 56700 12898 56756 12910
rect 56812 12962 57316 12964
rect 56812 12910 57262 12962
rect 57314 12910 57316 12962
rect 56812 12908 57316 12910
rect 56700 12404 56756 12414
rect 56700 12178 56756 12348
rect 56700 12126 56702 12178
rect 56754 12126 56756 12178
rect 56700 11956 56756 12126
rect 56700 11890 56756 11900
rect 56812 11732 56868 12908
rect 57260 12898 57316 12908
rect 57036 12738 57092 12750
rect 57036 12686 57038 12738
rect 57090 12686 57092 12738
rect 57036 12404 57092 12686
rect 57148 12740 57204 12750
rect 57148 12646 57204 12684
rect 57484 12738 57540 12750
rect 57484 12686 57486 12738
rect 57538 12686 57540 12738
rect 57484 12404 57540 12686
rect 57036 12348 57428 12404
rect 56588 11676 56868 11732
rect 57148 12178 57204 12190
rect 57148 12126 57150 12178
rect 57202 12126 57204 12178
rect 56140 10782 56142 10834
rect 56194 10782 56196 10834
rect 56140 10770 56196 10782
rect 56252 11394 56308 11406
rect 56252 11342 56254 11394
rect 56306 11342 56308 11394
rect 56252 10836 56308 11342
rect 56252 10770 56308 10780
rect 56364 11284 56420 11294
rect 56364 11170 56420 11228
rect 56364 11118 56366 11170
rect 56418 11118 56420 11170
rect 55580 10670 55582 10722
rect 55634 10670 55636 10722
rect 55580 10658 55636 10670
rect 56364 10612 56420 11118
rect 55020 6802 55076 7980
rect 55020 6750 55022 6802
rect 55074 6750 55076 6802
rect 55020 6738 55076 6750
rect 55244 10052 55300 10062
rect 55244 8930 55300 9996
rect 55356 9044 55412 9054
rect 55356 8950 55412 8988
rect 55244 8878 55246 8930
rect 55298 8878 55300 8930
rect 54908 6638 54910 6690
rect 54962 6638 54964 6690
rect 54908 6626 54964 6638
rect 54012 6078 54014 6130
rect 54066 6078 54068 6130
rect 54012 6066 54068 6078
rect 53900 5742 53902 5794
rect 53954 5742 53956 5794
rect 52220 5682 52276 5694
rect 52220 5630 52222 5682
rect 52274 5630 52276 5682
rect 51286 5516 51550 5526
rect 49532 5282 49588 5292
rect 50876 5460 50932 5470
rect 51342 5460 51390 5516
rect 51446 5460 51494 5516
rect 51286 5450 51550 5460
rect 49420 5236 49476 5246
rect 49308 5234 49476 5236
rect 49308 5182 49422 5234
rect 49474 5182 49476 5234
rect 49308 5180 49476 5182
rect 49420 5170 49476 5180
rect 49756 5236 49812 5246
rect 49756 5142 49812 5180
rect 50876 5234 50932 5404
rect 50876 5182 50878 5234
rect 50930 5182 50932 5234
rect 50876 5170 50932 5182
rect 51324 5348 51380 5358
rect 51324 5234 51380 5292
rect 51324 5182 51326 5234
rect 51378 5182 51380 5234
rect 51324 5170 51380 5182
rect 51100 5124 51156 5134
rect 49028 4844 49140 4900
rect 49644 4900 49700 4910
rect 48972 4562 49028 4844
rect 49644 4806 49700 4844
rect 49868 4900 49924 4910
rect 50428 4900 50484 4910
rect 49868 4898 50484 4900
rect 49868 4846 49870 4898
rect 49922 4846 50430 4898
rect 50482 4846 50484 4898
rect 49868 4844 50484 4846
rect 48972 4510 48974 4562
rect 49026 4510 49028 4562
rect 48972 4498 49028 4510
rect 49868 4564 49924 4844
rect 50428 4834 50484 4844
rect 49868 4498 49924 4508
rect 48524 3502 48526 3554
rect 48578 3502 48580 3554
rect 48524 3490 48580 3502
rect 48860 4452 48916 4462
rect 42700 3444 42756 3454
rect 42476 3442 42756 3444
rect 42476 3390 42702 3442
rect 42754 3390 42756 3442
rect 42476 3388 42756 3390
rect 48860 3444 48916 4396
rect 49308 4452 49364 4462
rect 49308 4338 49364 4396
rect 49308 4286 49310 4338
rect 49362 4286 49364 4338
rect 49308 4274 49364 4286
rect 49532 4338 49588 4350
rect 49532 4286 49534 4338
rect 49586 4286 49588 4338
rect 49532 4228 49588 4286
rect 51100 4338 51156 5068
rect 52220 5124 52276 5630
rect 53900 5460 53956 5742
rect 54012 5906 54068 5918
rect 54012 5854 54014 5906
rect 54066 5854 54068 5906
rect 54012 5796 54068 5854
rect 54012 5730 54068 5740
rect 54348 5906 54404 5918
rect 54348 5854 54350 5906
rect 54402 5854 54404 5906
rect 53900 5394 53956 5404
rect 54348 5348 54404 5854
rect 55244 5794 55300 8878
rect 55356 6692 55412 6702
rect 55468 6692 55524 10332
rect 56028 10556 56420 10612
rect 56028 9826 56084 10556
rect 56028 9774 56030 9826
rect 56082 9774 56084 9826
rect 56028 9762 56084 9774
rect 56476 9828 56532 9838
rect 56588 9828 56644 11676
rect 56700 11394 56756 11406
rect 56700 11342 56702 11394
rect 56754 11342 56756 11394
rect 56700 10052 56756 11342
rect 57148 11284 57204 12126
rect 57372 12178 57428 12348
rect 57484 12338 57540 12348
rect 57596 12402 57652 13694
rect 57596 12350 57598 12402
rect 57650 12350 57652 12402
rect 57596 12338 57652 12350
rect 57708 12292 57764 12302
rect 57708 12198 57764 12236
rect 57372 12126 57374 12178
rect 57426 12126 57428 12178
rect 57260 12066 57316 12078
rect 57260 12014 57262 12066
rect 57314 12014 57316 12066
rect 57260 11844 57316 12014
rect 57260 11778 57316 11788
rect 57148 11218 57204 11228
rect 57372 11172 57428 12126
rect 57820 12068 57876 15092
rect 58439 14140 58703 14150
rect 58495 14084 58543 14140
rect 58599 14084 58647 14140
rect 58439 14074 58703 14084
rect 58156 13634 58212 13646
rect 58156 13582 58158 13634
rect 58210 13582 58212 13634
rect 58044 13412 58100 13422
rect 58044 13186 58100 13356
rect 58044 13134 58046 13186
rect 58098 13134 58100 13186
rect 58044 13122 58100 13134
rect 57932 12852 57988 12862
rect 57932 12758 57988 12796
rect 58044 12738 58100 12750
rect 58044 12686 58046 12738
rect 58098 12686 58100 12738
rect 57932 12180 57988 12190
rect 57932 12086 57988 12124
rect 57484 12012 57876 12068
rect 57484 11506 57540 12012
rect 58044 11956 58100 12686
rect 58156 12404 58212 13582
rect 58439 12572 58703 12582
rect 58495 12516 58543 12572
rect 58599 12516 58647 12572
rect 58439 12506 58703 12516
rect 58156 12338 58212 12348
rect 58156 12178 58212 12190
rect 58156 12126 58158 12178
rect 58210 12126 58212 12178
rect 58156 12068 58212 12126
rect 58156 12002 58212 12012
rect 57596 11900 58100 11956
rect 57596 11844 57652 11900
rect 57596 11778 57652 11788
rect 57484 11454 57486 11506
rect 57538 11454 57540 11506
rect 57484 11442 57540 11454
rect 57820 11732 57876 11742
rect 57820 11282 57876 11676
rect 57820 11230 57822 11282
rect 57874 11230 57876 11282
rect 57820 11218 57876 11230
rect 57372 11078 57428 11116
rect 57596 11170 57652 11182
rect 57596 11118 57598 11170
rect 57650 11118 57652 11170
rect 56924 10612 56980 10622
rect 56924 10518 56980 10556
rect 56700 9986 56756 9996
rect 56476 9826 57092 9828
rect 56476 9774 56478 9826
rect 56530 9774 57092 9826
rect 56476 9772 57092 9774
rect 56476 9762 56532 9772
rect 56476 9042 56532 9054
rect 56476 8990 56478 9042
rect 56530 8990 56532 9042
rect 56476 8484 56532 8990
rect 57036 8708 57092 9772
rect 57372 9716 57428 9726
rect 57596 9716 57652 11118
rect 58439 11004 58703 11014
rect 58495 10948 58543 11004
rect 58599 10948 58647 11004
rect 58439 10938 58703 10948
rect 57932 10386 57988 10398
rect 57932 10334 57934 10386
rect 57986 10334 57988 10386
rect 57932 10164 57988 10334
rect 57932 10098 57988 10108
rect 58156 9716 58212 9726
rect 57596 9714 58212 9716
rect 57596 9662 58158 9714
rect 58210 9662 58212 9714
rect 57596 9660 58212 9662
rect 57372 9154 57428 9660
rect 57372 9102 57374 9154
rect 57426 9102 57428 9154
rect 57372 9090 57428 9102
rect 57596 9042 57652 9054
rect 57596 8990 57598 9042
rect 57650 8990 57652 9042
rect 57036 8652 57204 8708
rect 56476 8370 56532 8428
rect 56476 8318 56478 8370
rect 56530 8318 56532 8370
rect 56476 8306 56532 8318
rect 57148 8370 57204 8652
rect 57148 8318 57150 8370
rect 57202 8318 57204 8370
rect 57148 8306 57204 8318
rect 55356 6690 55524 6692
rect 55356 6638 55358 6690
rect 55410 6638 55524 6690
rect 55356 6636 55524 6638
rect 55580 8260 55636 8270
rect 55356 6626 55412 6636
rect 55244 5742 55246 5794
rect 55298 5742 55300 5794
rect 55244 5684 55300 5742
rect 55468 5796 55524 5806
rect 55468 5702 55524 5740
rect 55356 5684 55412 5694
rect 55244 5628 55356 5684
rect 55356 5618 55412 5628
rect 55580 5572 55636 8204
rect 57260 8258 57316 8270
rect 57260 8206 57262 8258
rect 57314 8206 57316 8258
rect 57036 7588 57092 7598
rect 56812 7362 56868 7374
rect 56812 7310 56814 7362
rect 56866 7310 56868 7362
rect 56140 6692 56196 6702
rect 56140 6130 56196 6636
rect 56140 6078 56142 6130
rect 56194 6078 56196 6130
rect 56140 6066 56196 6078
rect 55692 6020 55748 6030
rect 55692 5906 55748 5964
rect 55692 5854 55694 5906
rect 55746 5854 55748 5906
rect 55692 5842 55748 5854
rect 55468 5516 55636 5572
rect 55692 5572 55748 5582
rect 55748 5516 56084 5572
rect 54348 5282 54404 5292
rect 55356 5460 55412 5470
rect 52220 5058 52276 5068
rect 54572 5124 54628 5134
rect 54572 5030 54628 5068
rect 55356 4788 55412 5404
rect 55468 5234 55524 5516
rect 55692 5460 55748 5516
rect 55468 5182 55470 5234
rect 55522 5182 55524 5234
rect 55468 5170 55524 5182
rect 55580 5404 55748 5460
rect 55580 5122 55636 5404
rect 55804 5348 55860 5358
rect 55580 5070 55582 5122
rect 55634 5070 55636 5122
rect 55580 5058 55636 5070
rect 55692 5236 55748 5246
rect 55356 4732 55524 4788
rect 51548 4452 51604 4462
rect 51548 4358 51604 4396
rect 51100 4286 51102 4338
rect 51154 4286 51156 4338
rect 51100 4274 51156 4286
rect 55468 4338 55524 4732
rect 55468 4286 55470 4338
rect 55522 4286 55524 4338
rect 55468 4274 55524 4286
rect 49532 4162 49588 4172
rect 50204 4228 50260 4238
rect 50652 4228 50708 4238
rect 50204 4226 50708 4228
rect 50204 4174 50206 4226
rect 50258 4174 50654 4226
rect 50706 4174 50708 4226
rect 50204 4172 50708 4174
rect 50204 4162 50260 4172
rect 50652 4162 50708 4172
rect 51286 3948 51550 3958
rect 51342 3892 51390 3948
rect 51446 3892 51494 3948
rect 51286 3882 51550 3892
rect 55580 3556 55636 3566
rect 55692 3556 55748 5180
rect 55804 5124 55860 5292
rect 55804 4562 55860 5068
rect 55804 4510 55806 4562
rect 55858 4510 55860 4562
rect 55804 4498 55860 4510
rect 56028 5236 56084 5516
rect 56028 4562 56084 5180
rect 56812 5236 56868 7310
rect 57036 6690 57092 7532
rect 57148 7476 57204 7486
rect 57148 6916 57204 7420
rect 57148 6850 57204 6860
rect 57036 6638 57038 6690
rect 57090 6638 57092 6690
rect 56924 5908 56980 5918
rect 56924 5814 56980 5852
rect 57036 5684 57092 6638
rect 56028 4510 56030 4562
rect 56082 4510 56084 4562
rect 56028 4498 56084 4510
rect 56588 5124 56644 5134
rect 55916 4228 55972 4238
rect 55916 4134 55972 4172
rect 56588 3666 56644 5068
rect 56812 3778 56868 5180
rect 56924 5628 57092 5684
rect 57260 6020 57316 8206
rect 57596 7588 57652 8990
rect 57596 7522 57652 7532
rect 57708 8930 57764 8942
rect 57708 8878 57710 8930
rect 57762 8878 57764 8930
rect 57708 8258 57764 8878
rect 57708 8206 57710 8258
rect 57762 8206 57764 8258
rect 57596 7362 57652 7374
rect 57596 7310 57598 7362
rect 57650 7310 57652 7362
rect 57372 6692 57428 6702
rect 57372 6598 57428 6636
rect 56924 4452 56980 5628
rect 56924 4386 56980 4396
rect 57036 5460 57092 5470
rect 56812 3726 56814 3778
rect 56866 3726 56868 3778
rect 56812 3714 56868 3726
rect 57036 3778 57092 5404
rect 57036 3726 57038 3778
rect 57090 3726 57092 3778
rect 57036 3714 57092 3726
rect 56588 3614 56590 3666
rect 56642 3614 56644 3666
rect 56588 3602 56644 3614
rect 55580 3554 55748 3556
rect 55580 3502 55582 3554
rect 55634 3502 55748 3554
rect 55580 3500 55748 3502
rect 55580 3490 55636 3500
rect 48972 3444 49028 3454
rect 48860 3442 49028 3444
rect 48860 3390 48974 3442
rect 49026 3390 49028 3442
rect 48860 3388 49028 3390
rect 42700 3378 42756 3388
rect 48972 3378 49028 3388
rect 56252 3442 56308 3454
rect 56252 3390 56254 3442
rect 56306 3390 56308 3442
rect 1820 3266 1876 3276
rect 15518 3164 15782 3174
rect 15574 3108 15622 3164
rect 15678 3108 15726 3164
rect 15518 3098 15782 3108
rect 29825 3164 30089 3174
rect 29881 3108 29929 3164
rect 29985 3108 30033 3164
rect 29825 3098 30089 3108
rect 44132 3164 44396 3174
rect 44188 3108 44236 3164
rect 44292 3108 44340 3164
rect 44132 3098 44396 3108
rect 56252 2996 56308 3390
rect 57260 3444 57316 5964
rect 57596 5796 57652 7310
rect 57484 5124 57540 5134
rect 57484 5030 57540 5068
rect 57596 4338 57652 5740
rect 57708 5684 57764 8206
rect 58044 7476 58100 7486
rect 58044 7382 58100 7420
rect 57932 7250 57988 7262
rect 57932 7198 57934 7250
rect 57986 7198 57988 7250
rect 57820 5684 57876 5694
rect 57708 5628 57820 5684
rect 57708 5460 57764 5470
rect 57708 5122 57764 5404
rect 57708 5070 57710 5122
rect 57762 5070 57764 5122
rect 57708 5058 57764 5070
rect 57596 4286 57598 4338
rect 57650 4286 57652 4338
rect 57596 4274 57652 4286
rect 57820 4338 57876 5628
rect 57932 5124 57988 7198
rect 58044 5908 58100 5918
rect 58044 5814 58100 5852
rect 57932 5058 57988 5068
rect 58044 4564 58100 4574
rect 58156 4564 58212 9660
rect 58439 9436 58703 9446
rect 58495 9380 58543 9436
rect 58599 9380 58647 9436
rect 58439 9370 58703 9380
rect 58439 7868 58703 7878
rect 58495 7812 58543 7868
rect 58599 7812 58647 7868
rect 58439 7802 58703 7812
rect 58439 6300 58703 6310
rect 58495 6244 58543 6300
rect 58599 6244 58647 6300
rect 58439 6234 58703 6244
rect 58439 4732 58703 4742
rect 58495 4676 58543 4732
rect 58599 4676 58647 4732
rect 58439 4666 58703 4676
rect 58044 4562 58212 4564
rect 58044 4510 58046 4562
rect 58098 4510 58212 4562
rect 58044 4508 58212 4510
rect 58044 4498 58100 4508
rect 57820 4286 57822 4338
rect 57874 4286 57876 4338
rect 57820 4274 57876 4286
rect 57932 4228 57988 4238
rect 57484 3668 57540 3678
rect 57484 3666 57876 3668
rect 57484 3614 57486 3666
rect 57538 3614 57876 3666
rect 57484 3612 57876 3614
rect 57484 3602 57540 3612
rect 57596 3444 57652 3454
rect 57260 3442 57652 3444
rect 57260 3390 57598 3442
rect 57650 3390 57652 3442
rect 57260 3388 57652 3390
rect 57596 3378 57652 3388
rect 57820 3442 57876 3612
rect 57932 3554 57988 4172
rect 57932 3502 57934 3554
rect 57986 3502 57988 3554
rect 57932 3490 57988 3502
rect 57820 3390 57822 3442
rect 57874 3390 57876 3442
rect 57820 3378 57876 3390
rect 58439 3164 58703 3174
rect 58495 3108 58543 3164
rect 58599 3108 58647 3164
rect 58439 3098 58703 3108
rect 56252 2930 56308 2940
rect 1708 1362 1764 1372
<< via2 >>
rect 5516 28252 5572 28308
rect 2156 26460 2212 26516
rect 1484 26348 1540 26404
rect 1260 26012 1316 26068
rect 1260 13132 1316 13188
rect 1708 24668 1764 24724
rect 7980 26460 8036 26516
rect 4060 25676 4116 25732
rect 3052 25340 3108 25396
rect 2156 23436 2212 23492
rect 2268 23100 2324 23156
rect 1820 22764 1876 22820
rect 1708 21756 1764 21812
rect 4844 25228 4900 25284
rect 2940 23266 2996 23268
rect 2940 23214 2942 23266
rect 2942 23214 2994 23266
rect 2994 23214 2996 23266
rect 2940 23212 2996 23214
rect 2604 22876 2660 22932
rect 2716 22764 2772 22820
rect 1708 21084 1764 21140
rect 2604 21756 2660 21812
rect 1708 19292 1764 19348
rect 2268 20300 2324 20356
rect 2940 20300 2996 20356
rect 2716 20188 2772 20244
rect 2044 20018 2100 20020
rect 2044 19966 2046 20018
rect 2046 19966 2098 20018
rect 2098 19966 2100 20018
rect 2044 19964 2100 19966
rect 2492 19740 2548 19796
rect 1932 18284 1988 18340
rect 1820 17500 1876 17556
rect 1484 13020 1540 13076
rect 1596 15708 1652 15764
rect 2044 17724 2100 17780
rect 2828 18450 2884 18452
rect 2828 18398 2830 18450
rect 2830 18398 2882 18450
rect 2882 18398 2884 18450
rect 2828 18396 2884 18398
rect 2044 16770 2100 16772
rect 2044 16718 2046 16770
rect 2046 16718 2098 16770
rect 2098 16718 2100 16770
rect 2044 16716 2100 16718
rect 1932 15260 1988 15316
rect 1820 14812 1876 14868
rect 1820 14588 1876 14644
rect 1708 13916 1764 13972
rect 2268 17052 2324 17108
rect 2940 17778 2996 17780
rect 2940 17726 2942 17778
rect 2942 17726 2994 17778
rect 2994 17726 2996 17778
rect 2940 17724 2996 17726
rect 3276 24050 3332 24052
rect 3276 23998 3278 24050
rect 3278 23998 3330 24050
rect 3330 23998 3332 24050
rect 3276 23996 3332 23998
rect 4732 24668 4788 24724
rect 4620 23826 4676 23828
rect 4620 23774 4622 23826
rect 4622 23774 4674 23826
rect 4674 23774 4676 23826
rect 4620 23772 4676 23774
rect 3724 23212 3780 23268
rect 4732 23212 4788 23268
rect 3836 23100 3892 23156
rect 3388 21810 3444 21812
rect 3388 21758 3390 21810
rect 3390 21758 3442 21810
rect 3442 21758 3444 21810
rect 3388 21756 3444 21758
rect 3500 21586 3556 21588
rect 3500 21534 3502 21586
rect 3502 21534 3554 21586
rect 3554 21534 3556 21586
rect 3500 21532 3556 21534
rect 4620 23100 4676 23156
rect 4060 22876 4116 22932
rect 3276 20690 3332 20692
rect 3276 20638 3278 20690
rect 3278 20638 3330 20690
rect 3330 20638 3332 20690
rect 3276 20636 3332 20638
rect 3612 20300 3668 20356
rect 3164 20018 3220 20020
rect 3164 19966 3166 20018
rect 3166 19966 3218 20018
rect 3218 19966 3220 20018
rect 3164 19964 3220 19966
rect 2268 16828 2324 16884
rect 2268 16380 2324 16436
rect 3388 19964 3444 20020
rect 3500 19180 3556 19236
rect 3388 17164 3444 17220
rect 3052 17052 3108 17108
rect 2940 16716 2996 16772
rect 2716 16492 2772 16548
rect 2492 16268 2548 16324
rect 2268 15372 2324 15428
rect 3164 16380 3220 16436
rect 2604 15426 2660 15428
rect 2604 15374 2606 15426
rect 2606 15374 2658 15426
rect 2658 15374 2660 15426
rect 2604 15372 2660 15374
rect 2828 15372 2884 15428
rect 2716 15260 2772 15316
rect 2156 14812 2212 14868
rect 2604 15036 2660 15092
rect 2940 14530 2996 14532
rect 2940 14478 2942 14530
rect 2942 14478 2994 14530
rect 2994 14478 2996 14530
rect 2940 14476 2996 14478
rect 2268 14028 2324 14084
rect 1932 13634 1988 13636
rect 1932 13582 1934 13634
rect 1934 13582 1986 13634
rect 1986 13582 1988 13634
rect 1932 13580 1988 13582
rect 1932 12796 1988 12852
rect 2156 12796 2212 12852
rect 2156 12124 2212 12180
rect 2044 11340 2100 11396
rect 1932 10220 1988 10276
rect 1932 9660 1988 9716
rect 2716 13804 2772 13860
rect 2268 11900 2324 11956
rect 2380 13580 2436 13636
rect 3052 13468 3108 13524
rect 3164 14812 3220 14868
rect 2940 13356 2996 13412
rect 2380 11564 2436 11620
rect 2492 11676 2548 11732
rect 3164 12460 3220 12516
rect 2828 12012 2884 12068
rect 2940 11788 2996 11844
rect 3948 19852 4004 19908
rect 3948 18562 4004 18564
rect 3948 18510 3950 18562
rect 3950 18510 4002 18562
rect 4002 18510 4004 18562
rect 3948 18508 4004 18510
rect 3836 18450 3892 18452
rect 3836 18398 3838 18450
rect 3838 18398 3890 18450
rect 3890 18398 3892 18450
rect 3836 18396 3892 18398
rect 3612 17724 3668 17780
rect 3388 16156 3444 16212
rect 3500 16716 3556 16772
rect 3500 15372 3556 15428
rect 3724 16828 3780 16884
rect 3612 14140 3668 14196
rect 3500 13468 3556 13524
rect 3388 12124 3444 12180
rect 2268 10834 2324 10836
rect 2268 10782 2270 10834
rect 2270 10782 2322 10834
rect 2322 10782 2324 10834
rect 2268 10780 2324 10782
rect 3052 11340 3108 11396
rect 2940 10610 2996 10612
rect 2940 10558 2942 10610
rect 2942 10558 2994 10610
rect 2994 10558 2996 10610
rect 2940 10556 2996 10558
rect 3052 9772 3108 9828
rect 2492 8652 2548 8708
rect 2604 9660 2660 9716
rect 2380 8146 2436 8148
rect 2380 8094 2382 8146
rect 2382 8094 2434 8146
rect 2434 8094 2436 8146
rect 2380 8092 2436 8094
rect 1708 6690 1764 6692
rect 1708 6638 1710 6690
rect 1710 6638 1762 6690
rect 1762 6638 1764 6690
rect 1708 6636 1764 6638
rect 2492 7756 2548 7812
rect 2716 8540 2772 8596
rect 2716 8034 2772 8036
rect 2716 7982 2718 8034
rect 2718 7982 2770 8034
rect 2770 7982 2772 8034
rect 2716 7980 2772 7982
rect 3948 14364 4004 14420
rect 3836 13356 3892 13412
rect 3948 12684 4004 12740
rect 3948 12178 4004 12180
rect 3948 12126 3950 12178
rect 3950 12126 4002 12178
rect 4002 12126 4004 12178
rect 3948 12124 4004 12126
rect 3500 11170 3556 11172
rect 3500 11118 3502 11170
rect 3502 11118 3554 11170
rect 3554 11118 3556 11170
rect 3500 11116 3556 11118
rect 3388 9212 3444 9268
rect 3500 8988 3556 9044
rect 3612 9324 3668 9380
rect 3388 8876 3444 8932
rect 3948 11452 4004 11508
rect 3948 10892 4004 10948
rect 4284 19292 4340 19348
rect 5068 22988 5124 23044
rect 5180 23772 5236 23828
rect 4956 22876 5012 22932
rect 5404 23100 5460 23156
rect 5964 26178 6020 26180
rect 5964 26126 5966 26178
rect 5966 26126 6018 26178
rect 6018 26126 6020 26178
rect 5964 26124 6020 26126
rect 5852 25676 5908 25732
rect 7308 26290 7364 26292
rect 7308 26238 7310 26290
rect 7310 26238 7362 26290
rect 7362 26238 7364 26290
rect 7308 26236 7364 26238
rect 7196 25676 7252 25732
rect 7644 26012 7700 26068
rect 6860 25564 6916 25620
rect 7532 25564 7588 25620
rect 6972 25340 7028 25396
rect 5628 24834 5684 24836
rect 5628 24782 5630 24834
rect 5630 24782 5682 24834
rect 5682 24782 5684 24834
rect 5628 24780 5684 24782
rect 5628 22764 5684 22820
rect 4956 21868 5012 21924
rect 4396 18396 4452 18452
rect 4508 21532 4564 21588
rect 4508 20860 4564 20916
rect 4620 20748 4676 20804
rect 4732 20636 4788 20692
rect 4844 19906 4900 19908
rect 4844 19854 4846 19906
rect 4846 19854 4898 19906
rect 4898 19854 4900 19906
rect 4844 19852 4900 19854
rect 4508 17388 4564 17444
rect 4620 19122 4676 19124
rect 4620 19070 4622 19122
rect 4622 19070 4674 19122
rect 4674 19070 4676 19122
rect 4620 19068 4676 19070
rect 7196 25004 7252 25060
rect 7644 25228 7700 25284
rect 6636 24668 6692 24724
rect 6636 24498 6692 24500
rect 6636 24446 6638 24498
rect 6638 24446 6690 24498
rect 6690 24446 6692 24498
rect 6636 24444 6692 24446
rect 6412 23996 6468 24052
rect 6300 23042 6356 23044
rect 6300 22990 6302 23042
rect 6302 22990 6354 23042
rect 6354 22990 6356 23042
rect 6300 22988 6356 22990
rect 5180 21532 5236 21588
rect 6076 21586 6132 21588
rect 6076 21534 6078 21586
rect 6078 21534 6130 21586
rect 6130 21534 6132 21586
rect 6076 21532 6132 21534
rect 5964 21474 6020 21476
rect 5964 21422 5966 21474
rect 5966 21422 6018 21474
rect 6018 21422 6020 21474
rect 5964 21420 6020 21422
rect 5852 20860 5908 20916
rect 5180 20300 5236 20356
rect 5740 19068 5796 19124
rect 5068 19010 5124 19012
rect 5068 18958 5070 19010
rect 5070 18958 5122 19010
rect 5122 18958 5124 19010
rect 5068 18956 5124 18958
rect 4732 17442 4788 17444
rect 4732 17390 4734 17442
rect 4734 17390 4786 17442
rect 4786 17390 4788 17442
rect 4732 17388 4788 17390
rect 4620 16940 4676 16996
rect 4508 16828 4564 16884
rect 4172 16156 4228 16212
rect 4396 15426 4452 15428
rect 4396 15374 4398 15426
rect 4398 15374 4450 15426
rect 4450 15374 4452 15426
rect 4396 15372 4452 15374
rect 4732 15484 4788 15540
rect 5292 18620 5348 18676
rect 6076 19180 6132 19236
rect 5740 18562 5796 18564
rect 5740 18510 5742 18562
rect 5742 18510 5794 18562
rect 5794 18510 5796 18562
rect 5740 18508 5796 18510
rect 6076 18450 6132 18452
rect 6076 18398 6078 18450
rect 6078 18398 6130 18450
rect 6130 18398 6132 18450
rect 6076 18396 6132 18398
rect 5628 17724 5684 17780
rect 5292 16716 5348 16772
rect 5516 17388 5572 17444
rect 6076 17778 6132 17780
rect 6076 17726 6078 17778
rect 6078 17726 6130 17778
rect 6130 17726 6132 17778
rect 6076 17724 6132 17726
rect 5740 16940 5796 16996
rect 5292 16492 5348 16548
rect 4508 14924 4564 14980
rect 4172 14140 4228 14196
rect 4284 14530 4340 14532
rect 4284 14478 4286 14530
rect 4286 14478 4338 14530
rect 4338 14478 4340 14530
rect 4284 14476 4340 14478
rect 4284 13916 4340 13972
rect 4284 12962 4340 12964
rect 4284 12910 4286 12962
rect 4286 12910 4338 12962
rect 4338 12910 4340 12962
rect 4284 12908 4340 12910
rect 4172 11676 4228 11732
rect 5292 15426 5348 15428
rect 5292 15374 5294 15426
rect 5294 15374 5346 15426
rect 5346 15374 5348 15426
rect 5292 15372 5348 15374
rect 6076 16716 6132 16772
rect 6076 16210 6132 16212
rect 6076 16158 6078 16210
rect 6078 16158 6130 16210
rect 6130 16158 6132 16210
rect 6076 16156 6132 16158
rect 5516 14924 5572 14980
rect 4732 12908 4788 12964
rect 4844 12236 4900 12292
rect 4844 11900 4900 11956
rect 4060 10780 4116 10836
rect 4172 11340 4228 11396
rect 3948 10332 4004 10388
rect 3836 9324 3892 9380
rect 4620 10556 4676 10612
rect 3836 9154 3892 9156
rect 3836 9102 3838 9154
rect 3838 9102 3890 9154
rect 3890 9102 3892 9154
rect 3836 9100 3892 9102
rect 4060 9042 4116 9044
rect 4060 8990 4062 9042
rect 4062 8990 4114 9042
rect 4114 8990 4116 9042
rect 4060 8988 4116 8990
rect 2828 7644 2884 7700
rect 2828 7474 2884 7476
rect 2828 7422 2830 7474
rect 2830 7422 2882 7474
rect 2882 7422 2884 7474
rect 2828 7420 2884 7422
rect 3388 7756 3444 7812
rect 3052 7420 3108 7476
rect 2380 7084 2436 7140
rect 1932 6300 1988 6356
rect 1820 6130 1876 6132
rect 1820 6078 1822 6130
rect 1822 6078 1874 6130
rect 1874 6078 1876 6130
rect 1820 6076 1876 6078
rect 2044 5964 2100 6020
rect 1820 4956 1876 5012
rect 1820 4508 1876 4564
rect 2380 5794 2436 5796
rect 2380 5742 2382 5794
rect 2382 5742 2434 5794
rect 2434 5742 2436 5794
rect 2380 5740 2436 5742
rect 2716 6636 2772 6692
rect 2716 6300 2772 6356
rect 2604 5906 2660 5908
rect 2604 5854 2606 5906
rect 2606 5854 2658 5906
rect 2658 5854 2660 5906
rect 2604 5852 2660 5854
rect 1820 3612 1876 3668
rect 1708 3388 1764 3444
rect 3052 7084 3108 7140
rect 2940 5682 2996 5684
rect 2940 5630 2942 5682
rect 2942 5630 2994 5682
rect 2994 5630 2996 5682
rect 2940 5628 2996 5630
rect 3164 5740 3220 5796
rect 3500 6636 3556 6692
rect 3948 8764 4004 8820
rect 3836 8540 3892 8596
rect 3836 8316 3892 8372
rect 3948 8204 4004 8260
rect 3836 8092 3892 8148
rect 4060 7980 4116 8036
rect 3836 5964 3892 6020
rect 3724 5852 3780 5908
rect 3836 5794 3892 5796
rect 3836 5742 3838 5794
rect 3838 5742 3890 5794
rect 3890 5742 3892 5794
rect 3836 5740 3892 5742
rect 3724 5628 3780 5684
rect 3724 5122 3780 5124
rect 3724 5070 3726 5122
rect 3726 5070 3778 5122
rect 3778 5070 3780 5122
rect 3724 5068 3780 5070
rect 4508 9772 4564 9828
rect 5964 15036 6020 15092
rect 5628 14140 5684 14196
rect 5068 13692 5124 13748
rect 5964 13858 6020 13860
rect 5964 13806 5966 13858
rect 5966 13806 6018 13858
rect 6018 13806 6020 13858
rect 5964 13804 6020 13806
rect 6300 22204 6356 22260
rect 6636 23714 6692 23716
rect 6636 23662 6638 23714
rect 6638 23662 6690 23714
rect 6690 23662 6692 23714
rect 6636 23660 6692 23662
rect 7196 23996 7252 24052
rect 7196 23772 7252 23828
rect 7532 23436 7588 23492
rect 7308 22764 7364 22820
rect 6300 21420 6356 21476
rect 6300 20972 6356 21028
rect 6412 20860 6468 20916
rect 6748 20802 6804 20804
rect 6748 20750 6750 20802
rect 6750 20750 6802 20802
rect 6802 20750 6804 20802
rect 6748 20748 6804 20750
rect 6860 20690 6916 20692
rect 6860 20638 6862 20690
rect 6862 20638 6914 20690
rect 6914 20638 6916 20690
rect 6860 20636 6916 20638
rect 6860 20412 6916 20468
rect 6748 18562 6804 18564
rect 6748 18510 6750 18562
rect 6750 18510 6802 18562
rect 6802 18510 6804 18562
rect 6748 18508 6804 18510
rect 7084 19906 7140 19908
rect 7084 19854 7086 19906
rect 7086 19854 7138 19906
rect 7138 19854 7140 19906
rect 7084 19852 7140 19854
rect 7196 19068 7252 19124
rect 7084 18508 7140 18564
rect 6972 18450 7028 18452
rect 6972 18398 6974 18450
rect 6974 18398 7026 18450
rect 7026 18398 7028 18450
rect 6972 18396 7028 18398
rect 7084 18284 7140 18340
rect 7084 17724 7140 17780
rect 7196 17836 7252 17892
rect 7084 17052 7140 17108
rect 6524 16882 6580 16884
rect 6524 16830 6526 16882
rect 6526 16830 6578 16882
rect 6578 16830 6580 16882
rect 6524 16828 6580 16830
rect 7084 16882 7140 16884
rect 7084 16830 7086 16882
rect 7086 16830 7138 16882
rect 7138 16830 7140 16882
rect 7084 16828 7140 16830
rect 6524 16156 6580 16212
rect 6636 15426 6692 15428
rect 6636 15374 6638 15426
rect 6638 15374 6690 15426
rect 6690 15374 6692 15426
rect 6636 15372 6692 15374
rect 7084 15372 7140 15428
rect 6300 14924 6356 14980
rect 6188 14476 6244 14532
rect 6412 14364 6468 14420
rect 6188 13746 6244 13748
rect 6188 13694 6190 13746
rect 6190 13694 6242 13746
rect 6242 13694 6244 13746
rect 6188 13692 6244 13694
rect 6076 13356 6132 13412
rect 5964 13074 6020 13076
rect 5964 13022 5966 13074
rect 5966 13022 6018 13074
rect 6018 13022 6020 13074
rect 5964 13020 6020 13022
rect 7420 21698 7476 21700
rect 7420 21646 7422 21698
rect 7422 21646 7474 21698
rect 7474 21646 7476 21698
rect 7420 21644 7476 21646
rect 7756 24444 7812 24500
rect 8092 25452 8148 25508
rect 9324 26402 9380 26404
rect 9324 26350 9326 26402
rect 9326 26350 9378 26402
rect 9378 26350 9380 26402
rect 9324 26348 9380 26350
rect 57708 27356 57764 27412
rect 15518 26682 15574 26684
rect 15518 26630 15520 26682
rect 15520 26630 15572 26682
rect 15572 26630 15574 26682
rect 15518 26628 15574 26630
rect 15622 26682 15678 26684
rect 15622 26630 15624 26682
rect 15624 26630 15676 26682
rect 15676 26630 15678 26682
rect 15622 26628 15678 26630
rect 15726 26682 15782 26684
rect 15726 26630 15728 26682
rect 15728 26630 15780 26682
rect 15780 26630 15782 26682
rect 15726 26628 15782 26630
rect 9884 26348 9940 26404
rect 10220 26236 10276 26292
rect 8876 26178 8932 26180
rect 8876 26126 8878 26178
rect 8878 26126 8930 26178
rect 8930 26126 8932 26178
rect 8876 26124 8932 26126
rect 8365 25898 8421 25900
rect 8365 25846 8367 25898
rect 8367 25846 8419 25898
rect 8419 25846 8421 25898
rect 8365 25844 8421 25846
rect 8469 25898 8525 25900
rect 8469 25846 8471 25898
rect 8471 25846 8523 25898
rect 8523 25846 8525 25898
rect 8469 25844 8525 25846
rect 8573 25898 8629 25900
rect 8573 25846 8575 25898
rect 8575 25846 8627 25898
rect 8627 25846 8629 25898
rect 8573 25844 8629 25846
rect 8764 25788 8820 25844
rect 9772 25788 9828 25844
rect 9436 25564 9492 25620
rect 9884 25676 9940 25732
rect 9100 25394 9156 25396
rect 9100 25342 9102 25394
rect 9102 25342 9154 25394
rect 9154 25342 9156 25394
rect 9100 25340 9156 25342
rect 8365 24330 8421 24332
rect 8365 24278 8367 24330
rect 8367 24278 8419 24330
rect 8419 24278 8421 24330
rect 8365 24276 8421 24278
rect 8469 24330 8525 24332
rect 8469 24278 8471 24330
rect 8471 24278 8523 24330
rect 8523 24278 8525 24330
rect 8469 24276 8525 24278
rect 8573 24330 8629 24332
rect 8573 24278 8575 24330
rect 8575 24278 8627 24330
rect 8627 24278 8629 24330
rect 8573 24276 8629 24278
rect 8204 24108 8260 24164
rect 8316 23772 8372 23828
rect 8988 25004 9044 25060
rect 8876 24108 8932 24164
rect 8988 23884 9044 23940
rect 9772 25340 9828 25396
rect 9884 24610 9940 24612
rect 9884 24558 9886 24610
rect 9886 24558 9938 24610
rect 9938 24558 9940 24610
rect 9884 24556 9940 24558
rect 10220 24108 10276 24164
rect 8092 22428 8148 22484
rect 8365 22762 8421 22764
rect 8365 22710 8367 22762
rect 8367 22710 8419 22762
rect 8419 22710 8421 22762
rect 8365 22708 8421 22710
rect 8469 22762 8525 22764
rect 8469 22710 8471 22762
rect 8471 22710 8523 22762
rect 8523 22710 8525 22762
rect 8469 22708 8525 22710
rect 8573 22762 8629 22764
rect 8573 22710 8575 22762
rect 8575 22710 8627 22762
rect 8627 22710 8629 22762
rect 8573 22708 8629 22710
rect 9100 23100 9156 23156
rect 8876 22876 8932 22932
rect 8204 22258 8260 22260
rect 8204 22206 8206 22258
rect 8206 22206 8258 22258
rect 8258 22206 8260 22258
rect 8204 22204 8260 22206
rect 8876 22370 8932 22372
rect 8876 22318 8878 22370
rect 8878 22318 8930 22370
rect 8930 22318 8932 22370
rect 8876 22316 8932 22318
rect 8876 21810 8932 21812
rect 8876 21758 8878 21810
rect 8878 21758 8930 21810
rect 8930 21758 8932 21810
rect 8876 21756 8932 21758
rect 7756 20578 7812 20580
rect 7756 20526 7758 20578
rect 7758 20526 7810 20578
rect 7810 20526 7812 20578
rect 7756 20524 7812 20526
rect 7644 19964 7700 20020
rect 7644 18844 7700 18900
rect 7420 18508 7476 18564
rect 7420 15596 7476 15652
rect 6636 14476 6692 14532
rect 6748 14252 6804 14308
rect 6860 13970 6916 13972
rect 6860 13918 6862 13970
rect 6862 13918 6914 13970
rect 6914 13918 6916 13970
rect 6860 13916 6916 13918
rect 6972 13356 7028 13412
rect 5852 11788 5908 11844
rect 5740 11676 5796 11732
rect 5292 11116 5348 11172
rect 4956 10498 5012 10500
rect 4956 10446 4958 10498
rect 4958 10446 5010 10498
rect 5010 10446 5012 10498
rect 4956 10444 5012 10446
rect 4508 9436 4564 9492
rect 4844 9436 4900 9492
rect 4508 9154 4564 9156
rect 4508 9102 4510 9154
rect 4510 9102 4562 9154
rect 4562 9102 4564 9154
rect 4508 9100 4564 9102
rect 4844 9154 4900 9156
rect 4844 9102 4846 9154
rect 4846 9102 4898 9154
rect 4898 9102 4900 9154
rect 4844 9100 4900 9102
rect 5068 9324 5124 9380
rect 4956 8876 5012 8932
rect 4396 8764 4452 8820
rect 5180 8764 5236 8820
rect 4508 8428 4564 8484
rect 4844 8652 4900 8708
rect 4844 8370 4900 8372
rect 4844 8318 4846 8370
rect 4846 8318 4898 8370
rect 4898 8318 4900 8370
rect 4844 8316 4900 8318
rect 4396 7474 4452 7476
rect 4396 7422 4398 7474
rect 4398 7422 4450 7474
rect 4450 7422 4452 7474
rect 4396 7420 4452 7422
rect 4732 6802 4788 6804
rect 4732 6750 4734 6802
rect 4734 6750 4786 6802
rect 4786 6750 4788 6802
rect 4732 6748 4788 6750
rect 5516 10892 5572 10948
rect 5628 10610 5684 10612
rect 5628 10558 5630 10610
rect 5630 10558 5682 10610
rect 5682 10558 5684 10610
rect 5628 10556 5684 10558
rect 6300 11676 6356 11732
rect 6748 12348 6804 12404
rect 6188 11170 6244 11172
rect 6188 11118 6190 11170
rect 6190 11118 6242 11170
rect 6242 11118 6244 11170
rect 6188 11116 6244 11118
rect 6636 10556 6692 10612
rect 6076 9996 6132 10052
rect 7196 12738 7252 12740
rect 7196 12686 7198 12738
rect 7198 12686 7250 12738
rect 7250 12686 7252 12738
rect 7196 12684 7252 12686
rect 7308 11954 7364 11956
rect 7308 11902 7310 11954
rect 7310 11902 7362 11954
rect 7362 11902 7364 11954
rect 7308 11900 7364 11902
rect 6860 9996 6916 10052
rect 6300 9826 6356 9828
rect 6300 9774 6302 9826
rect 6302 9774 6354 9826
rect 6354 9774 6356 9826
rect 6300 9772 6356 9774
rect 6300 9212 6356 9268
rect 6748 9212 6804 9268
rect 8988 21586 9044 21588
rect 8988 21534 8990 21586
rect 8990 21534 9042 21586
rect 9042 21534 9044 21586
rect 8988 21532 9044 21534
rect 8365 21194 8421 21196
rect 8365 21142 8367 21194
rect 8367 21142 8419 21194
rect 8419 21142 8421 21194
rect 8365 21140 8421 21142
rect 8469 21194 8525 21196
rect 8469 21142 8471 21194
rect 8471 21142 8523 21194
rect 8523 21142 8525 21194
rect 8469 21140 8525 21142
rect 8573 21194 8629 21196
rect 8573 21142 8575 21194
rect 8575 21142 8627 21194
rect 8627 21142 8629 21194
rect 8573 21140 8629 21142
rect 9100 20412 9156 20468
rect 8428 20188 8484 20244
rect 8764 19852 8820 19908
rect 8365 19626 8421 19628
rect 8365 19574 8367 19626
rect 8367 19574 8419 19626
rect 8419 19574 8421 19626
rect 8365 19572 8421 19574
rect 8469 19626 8525 19628
rect 8469 19574 8471 19626
rect 8471 19574 8523 19626
rect 8523 19574 8525 19626
rect 8469 19572 8525 19574
rect 8573 19626 8629 19628
rect 8573 19574 8575 19626
rect 8575 19574 8627 19626
rect 8627 19574 8629 19626
rect 8573 19572 8629 19574
rect 8540 19122 8596 19124
rect 8540 19070 8542 19122
rect 8542 19070 8594 19122
rect 8594 19070 8596 19122
rect 8540 19068 8596 19070
rect 8876 19404 8932 19460
rect 9772 23154 9828 23156
rect 9772 23102 9774 23154
rect 9774 23102 9826 23154
rect 9826 23102 9828 23154
rect 9772 23100 9828 23102
rect 10332 23938 10388 23940
rect 10332 23886 10334 23938
rect 10334 23886 10386 23938
rect 10386 23886 10388 23938
rect 10332 23884 10388 23886
rect 10108 20412 10164 20468
rect 10108 20188 10164 20244
rect 9996 20130 10052 20132
rect 9996 20078 9998 20130
rect 9998 20078 10050 20130
rect 10050 20078 10052 20130
rect 9996 20076 10052 20078
rect 9884 19906 9940 19908
rect 9884 19854 9886 19906
rect 9886 19854 9938 19906
rect 9938 19854 9940 19906
rect 9884 19852 9940 19854
rect 9324 19234 9380 19236
rect 9324 19182 9326 19234
rect 9326 19182 9378 19234
rect 9378 19182 9380 19234
rect 9324 19180 9380 19182
rect 8204 18620 8260 18676
rect 7980 18226 8036 18228
rect 7980 18174 7982 18226
rect 7982 18174 8034 18226
rect 8034 18174 8036 18226
rect 7980 18172 8036 18174
rect 8365 18058 8421 18060
rect 8365 18006 8367 18058
rect 8367 18006 8419 18058
rect 8419 18006 8421 18058
rect 8365 18004 8421 18006
rect 8469 18058 8525 18060
rect 8469 18006 8471 18058
rect 8471 18006 8523 18058
rect 8523 18006 8525 18058
rect 8469 18004 8525 18006
rect 8573 18058 8629 18060
rect 8573 18006 8575 18058
rect 8575 18006 8627 18058
rect 8627 18006 8629 18058
rect 8573 18004 8629 18006
rect 8204 17836 8260 17892
rect 7980 17724 8036 17780
rect 8876 18620 8932 18676
rect 8316 17666 8372 17668
rect 8316 17614 8318 17666
rect 8318 17614 8370 17666
rect 8370 17614 8372 17666
rect 8316 17612 8372 17614
rect 7868 16940 7924 16996
rect 8092 17276 8148 17332
rect 7868 16716 7924 16772
rect 8764 16828 8820 16884
rect 8365 16490 8421 16492
rect 8365 16438 8367 16490
rect 8367 16438 8419 16490
rect 8419 16438 8421 16490
rect 8365 16436 8421 16438
rect 8469 16490 8525 16492
rect 8469 16438 8471 16490
rect 8471 16438 8523 16490
rect 8523 16438 8525 16490
rect 8469 16436 8525 16438
rect 8573 16490 8629 16492
rect 8573 16438 8575 16490
rect 8575 16438 8627 16490
rect 8627 16438 8629 16490
rect 8573 16436 8629 16438
rect 8092 16156 8148 16212
rect 8540 16098 8596 16100
rect 8540 16046 8542 16098
rect 8542 16046 8594 16098
rect 8594 16046 8596 16098
rect 8540 16044 8596 16046
rect 8365 14922 8421 14924
rect 8365 14870 8367 14922
rect 8367 14870 8419 14922
rect 8419 14870 8421 14922
rect 8365 14868 8421 14870
rect 8469 14922 8525 14924
rect 8469 14870 8471 14922
rect 8471 14870 8523 14922
rect 8523 14870 8525 14922
rect 8469 14868 8525 14870
rect 8573 14922 8629 14924
rect 8573 14870 8575 14922
rect 8575 14870 8627 14922
rect 8627 14870 8629 14922
rect 8573 14868 8629 14870
rect 9100 18508 9156 18564
rect 9100 17052 9156 17108
rect 8988 16828 9044 16884
rect 8988 15372 9044 15428
rect 8988 14754 9044 14756
rect 8988 14702 8990 14754
rect 8990 14702 9042 14754
rect 9042 14702 9044 14754
rect 8988 14700 9044 14702
rect 9660 18338 9716 18340
rect 9660 18286 9662 18338
rect 9662 18286 9714 18338
rect 9714 18286 9716 18338
rect 9660 18284 9716 18286
rect 9772 17276 9828 17332
rect 9660 16882 9716 16884
rect 9660 16830 9662 16882
rect 9662 16830 9714 16882
rect 9714 16830 9716 16882
rect 9660 16828 9716 16830
rect 9772 16716 9828 16772
rect 9660 15426 9716 15428
rect 9660 15374 9662 15426
rect 9662 15374 9714 15426
rect 9714 15374 9716 15426
rect 9660 15372 9716 15374
rect 10332 20524 10388 20580
rect 10220 19964 10276 20020
rect 10108 18956 10164 19012
rect 10220 19404 10276 19460
rect 11340 26290 11396 26292
rect 11340 26238 11342 26290
rect 11342 26238 11394 26290
rect 11394 26238 11396 26290
rect 11340 26236 11396 26238
rect 11116 26012 11172 26068
rect 12012 25618 12068 25620
rect 12012 25566 12014 25618
rect 12014 25566 12066 25618
rect 12066 25566 12068 25618
rect 12012 25564 12068 25566
rect 11452 25228 11508 25284
rect 11900 25452 11956 25508
rect 12460 25452 12516 25508
rect 12348 25282 12404 25284
rect 12348 25230 12350 25282
rect 12350 25230 12402 25282
rect 12402 25230 12404 25282
rect 12348 25228 12404 25230
rect 10892 24668 10948 24724
rect 10780 23660 10836 23716
rect 10556 21420 10612 21476
rect 11004 24108 11060 24164
rect 13580 26460 13636 26516
rect 13244 25564 13300 25620
rect 21308 26514 21364 26516
rect 21308 26462 21310 26514
rect 21310 26462 21362 26514
rect 21362 26462 21364 26514
rect 21308 26460 21364 26462
rect 26684 26460 26740 26516
rect 13468 25506 13524 25508
rect 13468 25454 13470 25506
rect 13470 25454 13522 25506
rect 13522 25454 13524 25506
rect 13468 25452 13524 25454
rect 12236 24668 12292 24724
rect 11900 23884 11956 23940
rect 12236 23996 12292 24052
rect 11676 23324 11732 23380
rect 11900 23100 11956 23156
rect 11452 21868 11508 21924
rect 10668 21644 10724 21700
rect 10556 20018 10612 20020
rect 10556 19966 10558 20018
rect 10558 19966 10610 20018
rect 10610 19966 10612 20018
rect 10556 19964 10612 19966
rect 10444 19180 10500 19236
rect 11564 21532 11620 21588
rect 10780 21420 10836 21476
rect 10892 20972 10948 21028
rect 10780 18956 10836 19012
rect 10220 18732 10276 18788
rect 10332 18844 10388 18900
rect 10780 18620 10836 18676
rect 10332 18508 10388 18564
rect 10668 18226 10724 18228
rect 10668 18174 10670 18226
rect 10670 18174 10722 18226
rect 10722 18174 10724 18226
rect 10668 18172 10724 18174
rect 10108 17500 10164 17556
rect 9996 16268 10052 16324
rect 10444 17388 10500 17444
rect 11676 21868 11732 21924
rect 12572 24668 12628 24724
rect 13356 24722 13412 24724
rect 13356 24670 13358 24722
rect 13358 24670 13410 24722
rect 13410 24670 13412 24722
rect 13356 24668 13412 24670
rect 12908 24050 12964 24052
rect 12908 23998 12910 24050
rect 12910 23998 12962 24050
rect 12962 23998 12964 24050
rect 12908 23996 12964 23998
rect 13356 23884 13412 23940
rect 13468 24556 13524 24612
rect 13468 24220 13524 24276
rect 12236 23548 12292 23604
rect 13132 23212 13188 23268
rect 12684 23154 12740 23156
rect 12684 23102 12686 23154
rect 12686 23102 12738 23154
rect 12738 23102 12740 23154
rect 12684 23100 12740 23102
rect 13020 21868 13076 21924
rect 11900 21420 11956 21476
rect 11452 20188 11508 20244
rect 11228 19964 11284 20020
rect 11116 19180 11172 19236
rect 11004 18284 11060 18340
rect 11004 17778 11060 17780
rect 11004 17726 11006 17778
rect 11006 17726 11058 17778
rect 11058 17726 11060 17778
rect 11004 17724 11060 17726
rect 11004 16994 11060 16996
rect 11004 16942 11006 16994
rect 11006 16942 11058 16994
rect 11058 16942 11060 16994
rect 11004 16940 11060 16942
rect 10892 16716 10948 16772
rect 10892 16380 10948 16436
rect 10556 15596 10612 15652
rect 11788 19180 11844 19236
rect 11564 18284 11620 18340
rect 11228 18060 11284 18116
rect 11004 15596 11060 15652
rect 9884 14700 9940 14756
rect 9996 14812 10052 14868
rect 8092 13580 8148 13636
rect 8204 14252 8260 14308
rect 9436 14306 9492 14308
rect 9436 14254 9438 14306
rect 9438 14254 9490 14306
rect 9490 14254 9492 14306
rect 9436 14252 9492 14254
rect 9772 14140 9828 14196
rect 9660 13634 9716 13636
rect 9660 13582 9662 13634
rect 9662 13582 9714 13634
rect 9714 13582 9716 13634
rect 9660 13580 9716 13582
rect 8764 13522 8820 13524
rect 8764 13470 8766 13522
rect 8766 13470 8818 13522
rect 8818 13470 8820 13522
rect 8764 13468 8820 13470
rect 8365 13354 8421 13356
rect 8365 13302 8367 13354
rect 8367 13302 8419 13354
rect 8419 13302 8421 13354
rect 8365 13300 8421 13302
rect 8469 13354 8525 13356
rect 8469 13302 8471 13354
rect 8471 13302 8523 13354
rect 8523 13302 8525 13354
rect 8469 13300 8525 13302
rect 8573 13354 8629 13356
rect 8573 13302 8575 13354
rect 8575 13302 8627 13354
rect 8627 13302 8629 13354
rect 8573 13300 8629 13302
rect 9436 12850 9492 12852
rect 9436 12798 9438 12850
rect 9438 12798 9490 12850
rect 9490 12798 9492 12850
rect 9436 12796 9492 12798
rect 9660 12402 9716 12404
rect 9660 12350 9662 12402
rect 9662 12350 9714 12402
rect 9714 12350 9716 12402
rect 9660 12348 9716 12350
rect 8988 12124 9044 12180
rect 7420 10610 7476 10612
rect 7420 10558 7422 10610
rect 7422 10558 7474 10610
rect 7474 10558 7476 10610
rect 7420 10556 7476 10558
rect 8365 11786 8421 11788
rect 8365 11734 8367 11786
rect 8367 11734 8419 11786
rect 8419 11734 8421 11786
rect 8365 11732 8421 11734
rect 8469 11786 8525 11788
rect 8469 11734 8471 11786
rect 8471 11734 8523 11786
rect 8523 11734 8525 11786
rect 8469 11732 8525 11734
rect 8573 11786 8629 11788
rect 8573 11734 8575 11786
rect 8575 11734 8627 11786
rect 8627 11734 8629 11786
rect 8573 11732 8629 11734
rect 8764 11788 8820 11844
rect 8204 11340 8260 11396
rect 7868 11004 7924 11060
rect 7756 9996 7812 10052
rect 7084 9772 7140 9828
rect 7532 9266 7588 9268
rect 7532 9214 7534 9266
rect 7534 9214 7586 9266
rect 7586 9214 7588 9266
rect 7532 9212 7588 9214
rect 6076 8988 6132 9044
rect 6524 8988 6580 9044
rect 5404 8540 5460 8596
rect 4844 6076 4900 6132
rect 4172 5740 4228 5796
rect 4172 4732 4228 4788
rect 4620 5068 4676 5124
rect 4396 4562 4452 4564
rect 4396 4510 4398 4562
rect 4398 4510 4450 4562
rect 4450 4510 4452 4562
rect 4396 4508 4452 4510
rect 5740 8370 5796 8372
rect 5740 8318 5742 8370
rect 5742 8318 5794 8370
rect 5794 8318 5796 8370
rect 5740 8316 5796 8318
rect 6300 8204 6356 8260
rect 6636 8876 6692 8932
rect 6860 8540 6916 8596
rect 7420 8258 7476 8260
rect 7420 8206 7422 8258
rect 7422 8206 7474 8258
rect 7474 8206 7476 8258
rect 7420 8204 7476 8206
rect 6748 8146 6804 8148
rect 6748 8094 6750 8146
rect 6750 8094 6802 8146
rect 6802 8094 6804 8146
rect 6748 8092 6804 8094
rect 7308 8146 7364 8148
rect 7308 8094 7310 8146
rect 7310 8094 7362 8146
rect 7362 8094 7364 8146
rect 7308 8092 7364 8094
rect 7644 8540 7700 8596
rect 7756 9100 7812 9156
rect 5628 7868 5684 7924
rect 6188 7474 6244 7476
rect 6188 7422 6190 7474
rect 6190 7422 6242 7474
rect 6242 7422 6244 7474
rect 6188 7420 6244 7422
rect 5516 6636 5572 6692
rect 5740 6690 5796 6692
rect 5740 6638 5742 6690
rect 5742 6638 5794 6690
rect 5794 6638 5796 6690
rect 5740 6636 5796 6638
rect 5516 6130 5572 6132
rect 5516 6078 5518 6130
rect 5518 6078 5570 6130
rect 5570 6078 5572 6130
rect 5516 6076 5572 6078
rect 5740 5852 5796 5908
rect 5068 5068 5124 5124
rect 4956 4732 5012 4788
rect 5180 4562 5236 4564
rect 5180 4510 5182 4562
rect 5182 4510 5234 4562
rect 5234 4510 5236 4562
rect 5180 4508 5236 4510
rect 7532 7756 7588 7812
rect 7420 6636 7476 6692
rect 6972 6524 7028 6580
rect 7756 7756 7812 7812
rect 8316 10780 8372 10836
rect 8204 10556 8260 10612
rect 8092 9602 8148 9604
rect 8092 9550 8094 9602
rect 8094 9550 8146 9602
rect 8146 9550 8148 9602
rect 8092 9548 8148 9550
rect 8365 10218 8421 10220
rect 8365 10166 8367 10218
rect 8367 10166 8419 10218
rect 8419 10166 8421 10218
rect 8365 10164 8421 10166
rect 8469 10218 8525 10220
rect 8469 10166 8471 10218
rect 8471 10166 8523 10218
rect 8523 10166 8525 10218
rect 8469 10164 8525 10166
rect 8573 10218 8629 10220
rect 8573 10166 8575 10218
rect 8575 10166 8627 10218
rect 8627 10166 8629 10218
rect 8573 10164 8629 10166
rect 9548 12012 9604 12068
rect 9436 11394 9492 11396
rect 9436 11342 9438 11394
rect 9438 11342 9490 11394
rect 9490 11342 9492 11394
rect 9436 11340 9492 11342
rect 9100 9996 9156 10052
rect 9660 11788 9716 11844
rect 12012 19068 12068 19124
rect 11900 17836 11956 17892
rect 12012 18284 12068 18340
rect 12460 18508 12516 18564
rect 12348 18172 12404 18228
rect 11788 17612 11844 17668
rect 11676 17388 11732 17444
rect 11004 14588 11060 14644
rect 10108 11788 10164 11844
rect 9772 11564 9828 11620
rect 8988 9100 9044 9156
rect 9100 9826 9156 9828
rect 9100 9774 9102 9826
rect 9102 9774 9154 9826
rect 9154 9774 9156 9826
rect 9100 9772 9156 9774
rect 8540 8930 8596 8932
rect 8540 8878 8542 8930
rect 8542 8878 8594 8930
rect 8594 8878 8596 8930
rect 8540 8876 8596 8878
rect 8365 8650 8421 8652
rect 8365 8598 8367 8650
rect 8367 8598 8419 8650
rect 8419 8598 8421 8650
rect 8365 8596 8421 8598
rect 8469 8650 8525 8652
rect 8469 8598 8471 8650
rect 8471 8598 8523 8650
rect 8523 8598 8525 8650
rect 8469 8596 8525 8598
rect 8573 8650 8629 8652
rect 8573 8598 8575 8650
rect 8575 8598 8627 8650
rect 8627 8598 8629 8650
rect 8573 8596 8629 8598
rect 8876 8540 8932 8596
rect 8204 8258 8260 8260
rect 8204 8206 8206 8258
rect 8206 8206 8258 8258
rect 8258 8206 8260 8258
rect 8204 8204 8260 8206
rect 7980 8092 8036 8148
rect 9212 8146 9268 8148
rect 9212 8094 9214 8146
rect 9214 8094 9266 8146
rect 9266 8094 9268 8146
rect 9212 8092 9268 8094
rect 8428 7698 8484 7700
rect 8428 7646 8430 7698
rect 8430 7646 8482 7698
rect 8482 7646 8484 7698
rect 8428 7644 8484 7646
rect 9660 10892 9716 10948
rect 10108 10556 10164 10612
rect 9884 9772 9940 9828
rect 10108 9436 10164 9492
rect 9660 9266 9716 9268
rect 9660 9214 9662 9266
rect 9662 9214 9714 9266
rect 9714 9214 9716 9266
rect 9660 9212 9716 9214
rect 9772 9324 9828 9380
rect 10332 13074 10388 13076
rect 10332 13022 10334 13074
rect 10334 13022 10386 13074
rect 10386 13022 10388 13074
rect 10332 13020 10388 13022
rect 10444 12348 10500 12404
rect 10780 13804 10836 13860
rect 10668 13634 10724 13636
rect 10668 13582 10670 13634
rect 10670 13582 10722 13634
rect 10722 13582 10724 13634
rect 10668 13580 10724 13582
rect 10780 13356 10836 13412
rect 12348 17276 12404 17332
rect 11676 15260 11732 15316
rect 11452 14812 11508 14868
rect 11452 14476 11508 14532
rect 11340 13356 11396 13412
rect 11116 13074 11172 13076
rect 11116 13022 11118 13074
rect 11118 13022 11170 13074
rect 11170 13022 11172 13074
rect 11116 13020 11172 13022
rect 11564 14364 11620 14420
rect 12348 16098 12404 16100
rect 12348 16046 12350 16098
rect 12350 16046 12402 16098
rect 12402 16046 12404 16098
rect 12348 16044 12404 16046
rect 12012 15372 12068 15428
rect 12348 15314 12404 15316
rect 12348 15262 12350 15314
rect 12350 15262 12402 15314
rect 12402 15262 12404 15314
rect 12348 15260 12404 15262
rect 12124 14476 12180 14532
rect 12124 13580 12180 13636
rect 10668 12124 10724 12180
rect 11004 12402 11060 12404
rect 11004 12350 11006 12402
rect 11006 12350 11058 12402
rect 11058 12350 11060 12402
rect 11004 12348 11060 12350
rect 12796 19964 12852 20020
rect 12908 17666 12964 17668
rect 12908 17614 12910 17666
rect 12910 17614 12962 17666
rect 12962 17614 12964 17666
rect 12908 17612 12964 17614
rect 13020 17164 13076 17220
rect 12908 17052 12964 17108
rect 12684 15260 12740 15316
rect 12684 13020 12740 13076
rect 11676 12348 11732 12404
rect 12236 12348 12292 12404
rect 11340 11564 11396 11620
rect 10220 10386 10276 10388
rect 10220 10334 10222 10386
rect 10222 10334 10274 10386
rect 10274 10334 10276 10386
rect 10220 10332 10276 10334
rect 9996 9042 10052 9044
rect 9996 8990 9998 9042
rect 9998 8990 10050 9042
rect 10050 8990 10052 9042
rect 9996 8988 10052 8990
rect 9660 8540 9716 8596
rect 9772 8258 9828 8260
rect 9772 8206 9774 8258
rect 9774 8206 9826 8258
rect 9826 8206 9828 8258
rect 9772 8204 9828 8206
rect 10556 10444 10612 10500
rect 10444 9826 10500 9828
rect 10444 9774 10446 9826
rect 10446 9774 10498 9826
rect 10498 9774 10500 9826
rect 10444 9772 10500 9774
rect 10220 7980 10276 8036
rect 8365 7082 8421 7084
rect 8365 7030 8367 7082
rect 8367 7030 8419 7082
rect 8419 7030 8421 7082
rect 8365 7028 8421 7030
rect 8469 7082 8525 7084
rect 8469 7030 8471 7082
rect 8471 7030 8523 7082
rect 8523 7030 8525 7082
rect 8469 7028 8525 7030
rect 8573 7082 8629 7084
rect 8573 7030 8575 7082
rect 8575 7030 8627 7082
rect 8627 7030 8629 7082
rect 8573 7028 8629 7030
rect 11788 11618 11844 11620
rect 11788 11566 11790 11618
rect 11790 11566 11842 11618
rect 11842 11566 11844 11618
rect 11788 11564 11844 11566
rect 11676 11170 11732 11172
rect 11676 11118 11678 11170
rect 11678 11118 11730 11170
rect 11730 11118 11732 11170
rect 11676 11116 11732 11118
rect 11788 10668 11844 10724
rect 12124 11788 12180 11844
rect 12684 11788 12740 11844
rect 12908 11564 12964 11620
rect 12572 11506 12628 11508
rect 12572 11454 12574 11506
rect 12574 11454 12626 11506
rect 12626 11454 12628 11506
rect 12572 11452 12628 11454
rect 13020 11506 13076 11508
rect 13020 11454 13022 11506
rect 13022 11454 13074 11506
rect 13074 11454 13076 11506
rect 13020 11452 13076 11454
rect 12124 10722 12180 10724
rect 12124 10670 12126 10722
rect 12126 10670 12178 10722
rect 12178 10670 12180 10722
rect 12124 10668 12180 10670
rect 12572 10722 12628 10724
rect 12572 10670 12574 10722
rect 12574 10670 12626 10722
rect 12626 10670 12628 10722
rect 12572 10668 12628 10670
rect 12012 10556 12068 10612
rect 10668 9324 10724 9380
rect 10668 9154 10724 9156
rect 10668 9102 10670 9154
rect 10670 9102 10722 9154
rect 10722 9102 10724 9154
rect 10668 9100 10724 9102
rect 11228 9154 11284 9156
rect 11228 9102 11230 9154
rect 11230 9102 11282 9154
rect 11282 9102 11284 9154
rect 11228 9100 11284 9102
rect 10556 8316 10612 8372
rect 10444 8258 10500 8260
rect 10444 8206 10446 8258
rect 10446 8206 10498 8258
rect 10498 8206 10500 8258
rect 10444 8204 10500 8206
rect 10556 8092 10612 8148
rect 7756 5852 7812 5908
rect 7868 5740 7924 5796
rect 7308 5234 7364 5236
rect 7308 5182 7310 5234
rect 7310 5182 7362 5234
rect 7362 5182 7364 5234
rect 7308 5180 7364 5182
rect 6188 5122 6244 5124
rect 6188 5070 6190 5122
rect 6190 5070 6242 5122
rect 6242 5070 6244 5122
rect 6188 5068 6244 5070
rect 6636 4956 6692 5012
rect 6076 4732 6132 4788
rect 5628 4562 5684 4564
rect 5628 4510 5630 4562
rect 5630 4510 5682 4562
rect 5682 4510 5684 4562
rect 5628 4508 5684 4510
rect 4732 4284 4788 4340
rect 6300 4338 6356 4340
rect 6300 4286 6302 4338
rect 6302 4286 6354 4338
rect 6354 4286 6356 4338
rect 6300 4284 6356 4286
rect 4732 3666 4788 3668
rect 4732 3614 4734 3666
rect 4734 3614 4786 3666
rect 4786 3614 4788 3666
rect 4732 3612 4788 3614
rect 7196 4508 7252 4564
rect 6860 4284 6916 4340
rect 7532 4338 7588 4340
rect 7532 4286 7534 4338
rect 7534 4286 7586 4338
rect 7586 4286 7588 4338
rect 7532 4284 7588 4286
rect 13020 10332 13076 10388
rect 12796 9884 12852 9940
rect 12572 9100 12628 9156
rect 12012 8988 12068 9044
rect 12908 8764 12964 8820
rect 11564 8204 11620 8260
rect 12460 8258 12516 8260
rect 12460 8206 12462 8258
rect 12462 8206 12514 8258
rect 12514 8206 12516 8258
rect 12460 8204 12516 8206
rect 11228 8092 11284 8148
rect 10892 7980 10948 8036
rect 13580 23548 13636 23604
rect 13692 22316 13748 22372
rect 13468 22204 13524 22260
rect 13692 22092 13748 22148
rect 16044 26402 16100 26404
rect 16044 26350 16046 26402
rect 16046 26350 16098 26402
rect 16098 26350 16100 26402
rect 16044 26348 16100 26350
rect 15036 26066 15092 26068
rect 15036 26014 15038 26066
rect 15038 26014 15090 26066
rect 15090 26014 15092 26066
rect 15036 26012 15092 26014
rect 14364 25564 14420 25620
rect 14476 25452 14532 25508
rect 13804 21868 13860 21924
rect 13804 21644 13860 21700
rect 13692 18450 13748 18452
rect 13692 18398 13694 18450
rect 13694 18398 13746 18450
rect 13746 18398 13748 18450
rect 13692 18396 13748 18398
rect 13468 16380 13524 16436
rect 13356 16044 13412 16100
rect 13580 15932 13636 15988
rect 13468 14588 13524 14644
rect 14028 24108 14084 24164
rect 13916 21586 13972 21588
rect 13916 21534 13918 21586
rect 13918 21534 13970 21586
rect 13970 21534 13972 21586
rect 13916 21532 13972 21534
rect 14028 23884 14084 23940
rect 14140 22540 14196 22596
rect 15148 25506 15204 25508
rect 15148 25454 15150 25506
rect 15150 25454 15202 25506
rect 15202 25454 15204 25506
rect 15148 25452 15204 25454
rect 15518 25114 15574 25116
rect 15518 25062 15520 25114
rect 15520 25062 15572 25114
rect 15572 25062 15574 25114
rect 15518 25060 15574 25062
rect 15622 25114 15678 25116
rect 15622 25062 15624 25114
rect 15624 25062 15676 25114
rect 15676 25062 15678 25114
rect 15622 25060 15678 25062
rect 15726 25114 15782 25116
rect 15726 25062 15728 25114
rect 15728 25062 15780 25114
rect 15780 25062 15782 25114
rect 15726 25060 15782 25062
rect 14476 23884 14532 23940
rect 14476 21756 14532 21812
rect 15148 24722 15204 24724
rect 15148 24670 15150 24722
rect 15150 24670 15202 24722
rect 15202 24670 15204 24722
rect 15148 24668 15204 24670
rect 16380 26402 16436 26404
rect 16380 26350 16382 26402
rect 16382 26350 16434 26402
rect 16434 26350 16436 26402
rect 16380 26348 16436 26350
rect 20748 26402 20804 26404
rect 20748 26350 20750 26402
rect 20750 26350 20802 26402
rect 20802 26350 20804 26402
rect 20748 26348 20804 26350
rect 21532 26348 21588 26404
rect 16268 26290 16324 26292
rect 16268 26238 16270 26290
rect 16270 26238 16322 26290
rect 16322 26238 16324 26290
rect 16268 26236 16324 26238
rect 17500 26290 17556 26292
rect 17500 26238 17502 26290
rect 17502 26238 17554 26290
rect 17554 26238 17556 26290
rect 17500 26236 17556 26238
rect 16268 25340 16324 25396
rect 16716 25394 16772 25396
rect 16716 25342 16718 25394
rect 16718 25342 16770 25394
rect 16770 25342 16772 25394
rect 16716 25340 16772 25342
rect 16492 25282 16548 25284
rect 16492 25230 16494 25282
rect 16494 25230 16546 25282
rect 16546 25230 16548 25282
rect 16492 25228 16548 25230
rect 16044 24668 16100 24724
rect 15708 24444 15764 24500
rect 15260 23660 15316 23716
rect 16156 24108 16212 24164
rect 16044 23772 16100 23828
rect 15518 23546 15574 23548
rect 15518 23494 15520 23546
rect 15520 23494 15572 23546
rect 15572 23494 15574 23546
rect 15518 23492 15574 23494
rect 15622 23546 15678 23548
rect 15622 23494 15624 23546
rect 15624 23494 15676 23546
rect 15676 23494 15678 23546
rect 15622 23492 15678 23494
rect 15726 23546 15782 23548
rect 15726 23494 15728 23546
rect 15728 23494 15780 23546
rect 15780 23494 15782 23546
rect 15726 23492 15782 23494
rect 15036 22540 15092 22596
rect 16044 22540 16100 22596
rect 16044 22316 16100 22372
rect 15518 21978 15574 21980
rect 15518 21926 15520 21978
rect 15520 21926 15572 21978
rect 15572 21926 15574 21978
rect 15518 21924 15574 21926
rect 15622 21978 15678 21980
rect 15622 21926 15624 21978
rect 15624 21926 15676 21978
rect 15676 21926 15678 21978
rect 15622 21924 15678 21926
rect 15726 21978 15782 21980
rect 15726 21926 15728 21978
rect 15728 21926 15780 21978
rect 15780 21926 15782 21978
rect 15726 21924 15782 21926
rect 15932 21420 15988 21476
rect 15260 20748 15316 20804
rect 15148 20076 15204 20132
rect 14140 18620 14196 18676
rect 13916 15820 13972 15876
rect 14140 15314 14196 15316
rect 14140 15262 14142 15314
rect 14142 15262 14194 15314
rect 14194 15262 14196 15314
rect 14140 15260 14196 15262
rect 14364 19068 14420 19124
rect 15148 19404 15204 19460
rect 14700 18562 14756 18564
rect 14700 18510 14702 18562
rect 14702 18510 14754 18562
rect 14754 18510 14756 18562
rect 14700 18508 14756 18510
rect 15036 17836 15092 17892
rect 15518 20410 15574 20412
rect 15518 20358 15520 20410
rect 15520 20358 15572 20410
rect 15572 20358 15574 20410
rect 15518 20356 15574 20358
rect 15622 20410 15678 20412
rect 15622 20358 15624 20410
rect 15624 20358 15676 20410
rect 15676 20358 15678 20410
rect 15622 20356 15678 20358
rect 15726 20410 15782 20412
rect 15726 20358 15728 20410
rect 15728 20358 15780 20410
rect 15780 20358 15782 20410
rect 15726 20356 15782 20358
rect 15484 20076 15540 20132
rect 15820 20076 15876 20132
rect 15484 19628 15540 19684
rect 15596 20018 15652 20020
rect 15596 19966 15598 20018
rect 15598 19966 15650 20018
rect 15650 19966 15652 20018
rect 15596 19964 15652 19966
rect 16044 21362 16100 21364
rect 16044 21310 16046 21362
rect 16046 21310 16098 21362
rect 16098 21310 16100 21362
rect 16044 21308 16100 21310
rect 16044 20636 16100 20692
rect 15708 19234 15764 19236
rect 15708 19182 15710 19234
rect 15710 19182 15762 19234
rect 15762 19182 15764 19234
rect 15708 19180 15764 19182
rect 15260 18732 15316 18788
rect 15518 18842 15574 18844
rect 15518 18790 15520 18842
rect 15520 18790 15572 18842
rect 15572 18790 15574 18842
rect 15518 18788 15574 18790
rect 15622 18842 15678 18844
rect 15622 18790 15624 18842
rect 15624 18790 15676 18842
rect 15676 18790 15678 18842
rect 15622 18788 15678 18790
rect 15726 18842 15782 18844
rect 15726 18790 15728 18842
rect 15728 18790 15780 18842
rect 15780 18790 15782 18842
rect 15726 18788 15782 18790
rect 15484 18620 15540 18676
rect 15260 18508 15316 18564
rect 14364 17164 14420 17220
rect 14588 17052 14644 17108
rect 14476 15986 14532 15988
rect 14476 15934 14478 15986
rect 14478 15934 14530 15986
rect 14530 15934 14532 15986
rect 14476 15932 14532 15934
rect 15036 15874 15092 15876
rect 15036 15822 15038 15874
rect 15038 15822 15090 15874
rect 15090 15822 15092 15874
rect 15036 15820 15092 15822
rect 14924 15260 14980 15316
rect 13804 14588 13860 14644
rect 13580 12348 13636 12404
rect 14252 14812 14308 14868
rect 14252 14418 14308 14420
rect 14252 14366 14254 14418
rect 14254 14366 14306 14418
rect 14306 14366 14308 14418
rect 14252 14364 14308 14366
rect 14700 13244 14756 13300
rect 14364 12348 14420 12404
rect 13692 11506 13748 11508
rect 13692 11454 13694 11506
rect 13694 11454 13746 11506
rect 13746 11454 13748 11506
rect 13692 11452 13748 11454
rect 13580 11116 13636 11172
rect 13356 10556 13412 10612
rect 14140 11506 14196 11508
rect 14140 11454 14142 11506
rect 14142 11454 14194 11506
rect 14194 11454 14196 11506
rect 14140 11452 14196 11454
rect 15036 13858 15092 13860
rect 15036 13806 15038 13858
rect 15038 13806 15090 13858
rect 15090 13806 15092 13858
rect 15036 13804 15092 13806
rect 15148 15372 15204 15428
rect 15036 13244 15092 13300
rect 14588 11788 14644 11844
rect 14812 11900 14868 11956
rect 14140 11116 14196 11172
rect 14364 11116 14420 11172
rect 13692 9938 13748 9940
rect 13692 9886 13694 9938
rect 13694 9886 13746 9938
rect 13746 9886 13748 9938
rect 13692 9884 13748 9886
rect 13356 8764 13412 8820
rect 13580 8204 13636 8260
rect 14364 10444 14420 10500
rect 14700 10610 14756 10612
rect 14700 10558 14702 10610
rect 14702 10558 14754 10610
rect 14754 10558 14756 10610
rect 14700 10556 14756 10558
rect 14588 10332 14644 10388
rect 14252 9938 14308 9940
rect 14252 9886 14254 9938
rect 14254 9886 14306 9938
rect 14306 9886 14308 9938
rect 14252 9884 14308 9886
rect 13804 9772 13860 9828
rect 14476 9772 14532 9828
rect 13804 9154 13860 9156
rect 13804 9102 13806 9154
rect 13806 9102 13858 9154
rect 13858 9102 13860 9154
rect 13804 9100 13860 9102
rect 14700 9324 14756 9380
rect 14476 8764 14532 8820
rect 13132 7868 13188 7924
rect 12908 7644 12964 7700
rect 12124 7586 12180 7588
rect 12124 7534 12126 7586
rect 12126 7534 12178 7586
rect 12178 7534 12180 7586
rect 12124 7532 12180 7534
rect 11228 7474 11284 7476
rect 11228 7422 11230 7474
rect 11230 7422 11282 7474
rect 11282 7422 11284 7474
rect 11228 7420 11284 7422
rect 11900 7474 11956 7476
rect 11900 7422 11902 7474
rect 11902 7422 11954 7474
rect 11954 7422 11956 7474
rect 11900 7420 11956 7422
rect 13804 7644 13860 7700
rect 13916 7532 13972 7588
rect 14140 7420 14196 7476
rect 9996 6076 10052 6132
rect 8092 5180 8148 5236
rect 8316 5906 8372 5908
rect 8316 5854 8318 5906
rect 8318 5854 8370 5906
rect 8370 5854 8372 5906
rect 8316 5852 8372 5854
rect 8764 5906 8820 5908
rect 8764 5854 8766 5906
rect 8766 5854 8818 5906
rect 8818 5854 8820 5906
rect 8764 5852 8820 5854
rect 10108 5740 10164 5796
rect 8365 5514 8421 5516
rect 8365 5462 8367 5514
rect 8367 5462 8419 5514
rect 8419 5462 8421 5514
rect 8365 5460 8421 5462
rect 8469 5514 8525 5516
rect 8469 5462 8471 5514
rect 8471 5462 8523 5514
rect 8523 5462 8525 5514
rect 8469 5460 8525 5462
rect 8573 5514 8629 5516
rect 8573 5462 8575 5514
rect 8575 5462 8627 5514
rect 8627 5462 8629 5514
rect 8573 5460 8629 5462
rect 8316 5122 8372 5124
rect 8316 5070 8318 5122
rect 8318 5070 8370 5122
rect 8370 5070 8372 5122
rect 8316 5068 8372 5070
rect 9548 5010 9604 5012
rect 9548 4958 9550 5010
rect 9550 4958 9602 5010
rect 9602 4958 9604 5010
rect 9548 4956 9604 4958
rect 9772 4562 9828 4564
rect 9772 4510 9774 4562
rect 9774 4510 9826 4562
rect 9826 4510 9828 4562
rect 9772 4508 9828 4510
rect 8204 4450 8260 4452
rect 8204 4398 8206 4450
rect 8206 4398 8258 4450
rect 8258 4398 8260 4450
rect 8204 4396 8260 4398
rect 10220 5180 10276 5236
rect 10668 5740 10724 5796
rect 10780 5234 10836 5236
rect 10780 5182 10782 5234
rect 10782 5182 10834 5234
rect 10834 5182 10836 5234
rect 10780 5180 10836 5182
rect 10892 5122 10948 5124
rect 10892 5070 10894 5122
rect 10894 5070 10946 5122
rect 10946 5070 10948 5122
rect 10892 5068 10948 5070
rect 10668 4284 10724 4340
rect 12684 5852 12740 5908
rect 11676 5346 11732 5348
rect 11676 5294 11678 5346
rect 11678 5294 11730 5346
rect 11730 5294 11732 5346
rect 11676 5292 11732 5294
rect 12684 5292 12740 5348
rect 11004 4508 11060 4564
rect 11788 5180 11844 5236
rect 14588 7084 14644 7140
rect 14924 11788 14980 11844
rect 15260 14476 15316 14532
rect 16268 22316 16324 22372
rect 16268 22092 16324 22148
rect 16268 21308 16324 21364
rect 16828 24332 16884 24388
rect 16604 22092 16660 22148
rect 16716 23324 16772 23380
rect 16604 21756 16660 21812
rect 16716 20636 16772 20692
rect 16716 20412 16772 20468
rect 17276 23884 17332 23940
rect 16940 23378 16996 23380
rect 16940 23326 16942 23378
rect 16942 23326 16994 23378
rect 16994 23326 16996 23378
rect 16940 23324 16996 23326
rect 16940 22540 16996 22596
rect 17612 25506 17668 25508
rect 17612 25454 17614 25506
rect 17614 25454 17666 25506
rect 17666 25454 17668 25506
rect 17612 25452 17668 25454
rect 19628 26178 19684 26180
rect 19628 26126 19630 26178
rect 19630 26126 19682 26178
rect 19682 26126 19684 26178
rect 19628 26124 19684 26126
rect 19180 26012 19236 26068
rect 19964 26012 20020 26068
rect 19068 25452 19124 25508
rect 18732 25340 18788 25396
rect 18060 25228 18116 25284
rect 17500 24498 17556 24500
rect 17500 24446 17502 24498
rect 17502 24446 17554 24498
rect 17554 24446 17556 24498
rect 17500 24444 17556 24446
rect 17948 23884 18004 23940
rect 16940 21308 16996 21364
rect 17052 20802 17108 20804
rect 17052 20750 17054 20802
rect 17054 20750 17106 20802
rect 17106 20750 17108 20802
rect 17052 20748 17108 20750
rect 16492 20076 16548 20132
rect 16716 20076 16772 20132
rect 16156 19404 16212 19460
rect 16492 19516 16548 19572
rect 15820 18172 15876 18228
rect 16156 18226 16212 18228
rect 16156 18174 16158 18226
rect 16158 18174 16210 18226
rect 16210 18174 16212 18226
rect 16156 18172 16212 18174
rect 15518 17274 15574 17276
rect 15518 17222 15520 17274
rect 15520 17222 15572 17274
rect 15572 17222 15574 17274
rect 15518 17220 15574 17222
rect 15622 17274 15678 17276
rect 15622 17222 15624 17274
rect 15624 17222 15676 17274
rect 15676 17222 15678 17274
rect 15622 17220 15678 17222
rect 15726 17274 15782 17276
rect 15726 17222 15728 17274
rect 15728 17222 15780 17274
rect 15780 17222 15782 17274
rect 15726 17220 15782 17222
rect 16604 18620 16660 18676
rect 16492 18508 16548 18564
rect 15596 16994 15652 16996
rect 15596 16942 15598 16994
rect 15598 16942 15650 16994
rect 15650 16942 15652 16994
rect 15596 16940 15652 16942
rect 16828 18396 16884 18452
rect 15518 15706 15574 15708
rect 15518 15654 15520 15706
rect 15520 15654 15572 15706
rect 15572 15654 15574 15706
rect 15518 15652 15574 15654
rect 15622 15706 15678 15708
rect 15622 15654 15624 15706
rect 15624 15654 15676 15706
rect 15676 15654 15678 15706
rect 15622 15652 15678 15654
rect 15726 15706 15782 15708
rect 15726 15654 15728 15706
rect 15728 15654 15780 15706
rect 15780 15654 15782 15706
rect 15726 15652 15782 15654
rect 15484 15426 15540 15428
rect 15484 15374 15486 15426
rect 15486 15374 15538 15426
rect 15538 15374 15540 15426
rect 15484 15372 15540 15374
rect 16604 16658 16660 16660
rect 16604 16606 16606 16658
rect 16606 16606 16658 16658
rect 16658 16606 16660 16658
rect 16604 16604 16660 16606
rect 16268 15372 16324 15428
rect 16380 15314 16436 15316
rect 16380 15262 16382 15314
rect 16382 15262 16434 15314
rect 16434 15262 16436 15314
rect 16380 15260 16436 15262
rect 16156 15148 16212 15204
rect 16044 14530 16100 14532
rect 16044 14478 16046 14530
rect 16046 14478 16098 14530
rect 16098 14478 16100 14530
rect 16044 14476 16100 14478
rect 16044 14252 16100 14308
rect 15518 14138 15574 14140
rect 15518 14086 15520 14138
rect 15520 14086 15572 14138
rect 15572 14086 15574 14138
rect 15518 14084 15574 14086
rect 15622 14138 15678 14140
rect 15622 14086 15624 14138
rect 15624 14086 15676 14138
rect 15676 14086 15678 14138
rect 15622 14084 15678 14086
rect 15726 14138 15782 14140
rect 15726 14086 15728 14138
rect 15728 14086 15780 14138
rect 15780 14086 15782 14138
rect 15726 14084 15782 14086
rect 15708 13970 15764 13972
rect 15708 13918 15710 13970
rect 15710 13918 15762 13970
rect 15762 13918 15764 13970
rect 15708 13916 15764 13918
rect 15596 13804 15652 13860
rect 15372 13522 15428 13524
rect 15372 13470 15374 13522
rect 15374 13470 15426 13522
rect 15426 13470 15428 13522
rect 15372 13468 15428 13470
rect 16604 14364 16660 14420
rect 17836 23042 17892 23044
rect 17836 22990 17838 23042
rect 17838 22990 17890 23042
rect 17890 22990 17892 23042
rect 17836 22988 17892 22990
rect 17836 22540 17892 22596
rect 18396 24722 18452 24724
rect 18396 24670 18398 24722
rect 18398 24670 18450 24722
rect 18450 24670 18452 24722
rect 18396 24668 18452 24670
rect 18060 23212 18116 23268
rect 18508 24220 18564 24276
rect 18396 23548 18452 23604
rect 18284 22988 18340 23044
rect 18172 22092 18228 22148
rect 17612 21420 17668 21476
rect 17612 19964 17668 20020
rect 17052 19234 17108 19236
rect 17052 19182 17054 19234
rect 17054 19182 17106 19234
rect 17106 19182 17108 19234
rect 17052 19180 17108 19182
rect 17276 19628 17332 19684
rect 16940 18284 16996 18340
rect 17500 19404 17556 19460
rect 17388 18450 17444 18452
rect 17388 18398 17390 18450
rect 17390 18398 17442 18450
rect 17442 18398 17444 18450
rect 17388 18396 17444 18398
rect 17500 17724 17556 17780
rect 18620 22876 18676 22932
rect 18396 21980 18452 22036
rect 18284 18508 18340 18564
rect 18508 18844 18564 18900
rect 17724 18284 17780 18340
rect 16940 14812 16996 14868
rect 17164 16604 17220 16660
rect 18172 17666 18228 17668
rect 18172 17614 18174 17666
rect 18174 17614 18226 17666
rect 18226 17614 18228 17666
rect 18172 17612 18228 17614
rect 18396 17388 18452 17444
rect 19740 25340 19796 25396
rect 21084 26124 21140 26180
rect 20076 25788 20132 25844
rect 20972 25340 21028 25396
rect 20412 24332 20468 24388
rect 20636 24668 20692 24724
rect 19964 23938 20020 23940
rect 19964 23886 19966 23938
rect 19966 23886 20018 23938
rect 20018 23886 20020 23938
rect 19964 23884 20020 23886
rect 20076 24050 20132 24052
rect 20076 23998 20078 24050
rect 20078 23998 20130 24050
rect 20130 23998 20132 24050
rect 20076 23996 20132 23998
rect 20188 23324 20244 23380
rect 19628 22652 19684 22708
rect 19404 19852 19460 19908
rect 18844 18396 18900 18452
rect 19292 18508 19348 18564
rect 18732 18284 18788 18340
rect 19628 19010 19684 19012
rect 19628 18958 19630 19010
rect 19630 18958 19682 19010
rect 19682 18958 19684 19010
rect 19628 18956 19684 18958
rect 19740 18844 19796 18900
rect 18732 16828 18788 16884
rect 17724 15148 17780 15204
rect 17164 14418 17220 14420
rect 17164 14366 17166 14418
rect 17166 14366 17218 14418
rect 17218 14366 17220 14418
rect 17164 14364 17220 14366
rect 16716 14252 16772 14308
rect 16604 14028 16660 14084
rect 16940 14028 16996 14084
rect 16492 13916 16548 13972
rect 16716 13858 16772 13860
rect 16716 13806 16718 13858
rect 16718 13806 16770 13858
rect 16770 13806 16772 13858
rect 16716 13804 16772 13806
rect 16492 13468 16548 13524
rect 15518 12570 15574 12572
rect 15518 12518 15520 12570
rect 15520 12518 15572 12570
rect 15572 12518 15574 12570
rect 15518 12516 15574 12518
rect 15622 12570 15678 12572
rect 15622 12518 15624 12570
rect 15624 12518 15676 12570
rect 15676 12518 15678 12570
rect 15622 12516 15678 12518
rect 15726 12570 15782 12572
rect 15726 12518 15728 12570
rect 15728 12518 15780 12570
rect 15780 12518 15782 12570
rect 15726 12516 15782 12518
rect 16604 12908 16660 12964
rect 15260 11452 15316 11508
rect 15372 11564 15428 11620
rect 16380 12402 16436 12404
rect 16380 12350 16382 12402
rect 16382 12350 16434 12402
rect 16434 12350 16436 12402
rect 16380 12348 16436 12350
rect 17388 13970 17444 13972
rect 17388 13918 17390 13970
rect 17390 13918 17442 13970
rect 17442 13918 17444 13970
rect 17388 13916 17444 13918
rect 17612 13804 17668 13860
rect 18060 15932 18116 15988
rect 19404 17276 19460 17332
rect 19292 16882 19348 16884
rect 19292 16830 19294 16882
rect 19294 16830 19346 16882
rect 19346 16830 19348 16882
rect 19292 16828 19348 16830
rect 18844 16044 18900 16100
rect 18172 14812 18228 14868
rect 17948 13692 18004 13748
rect 16940 11900 16996 11956
rect 17052 13020 17108 13076
rect 16156 11564 16212 11620
rect 15260 10892 15316 10948
rect 15518 11002 15574 11004
rect 15518 10950 15520 11002
rect 15520 10950 15572 11002
rect 15572 10950 15574 11002
rect 15518 10948 15574 10950
rect 15622 11002 15678 11004
rect 15622 10950 15624 11002
rect 15624 10950 15676 11002
rect 15676 10950 15678 11002
rect 15622 10948 15678 10950
rect 15726 11002 15782 11004
rect 15726 10950 15728 11002
rect 15728 10950 15780 11002
rect 15780 10950 15782 11002
rect 15726 10948 15782 10950
rect 15148 10668 15204 10724
rect 15036 10556 15092 10612
rect 16604 10722 16660 10724
rect 16604 10670 16606 10722
rect 16606 10670 16658 10722
rect 16658 10670 16660 10722
rect 16604 10668 16660 10670
rect 15484 10556 15540 10612
rect 15372 10444 15428 10500
rect 15036 10332 15092 10388
rect 16268 10610 16324 10612
rect 16268 10558 16270 10610
rect 16270 10558 16322 10610
rect 16322 10558 16324 10610
rect 16268 10556 16324 10558
rect 16044 10386 16100 10388
rect 16044 10334 16046 10386
rect 16046 10334 16098 10386
rect 16098 10334 16100 10386
rect 16044 10332 16100 10334
rect 15708 9826 15764 9828
rect 15708 9774 15710 9826
rect 15710 9774 15762 9826
rect 15762 9774 15764 9826
rect 15708 9772 15764 9774
rect 15518 9434 15574 9436
rect 15518 9382 15520 9434
rect 15520 9382 15572 9434
rect 15572 9382 15574 9434
rect 15518 9380 15574 9382
rect 15622 9434 15678 9436
rect 15622 9382 15624 9434
rect 15624 9382 15676 9434
rect 15676 9382 15678 9434
rect 15622 9380 15678 9382
rect 15726 9434 15782 9436
rect 15726 9382 15728 9434
rect 15728 9382 15780 9434
rect 15780 9382 15782 9434
rect 15726 9380 15782 9382
rect 15596 9154 15652 9156
rect 15596 9102 15598 9154
rect 15598 9102 15650 9154
rect 15650 9102 15652 9154
rect 15596 9100 15652 9102
rect 14924 8764 14980 8820
rect 14924 8092 14980 8148
rect 15484 8540 15540 8596
rect 16156 9826 16212 9828
rect 16156 9774 16158 9826
rect 16158 9774 16210 9826
rect 16210 9774 16212 9826
rect 16156 9772 16212 9774
rect 17388 12908 17444 12964
rect 18620 14812 18676 14868
rect 18284 13916 18340 13972
rect 18396 14364 18452 14420
rect 18396 13804 18452 13860
rect 18172 12796 18228 12852
rect 17612 12066 17668 12068
rect 17612 12014 17614 12066
rect 17614 12014 17666 12066
rect 17666 12014 17668 12066
rect 17612 12012 17668 12014
rect 17500 11116 17556 11172
rect 17388 10722 17444 10724
rect 17388 10670 17390 10722
rect 17390 10670 17442 10722
rect 17442 10670 17444 10722
rect 17388 10668 17444 10670
rect 18284 12236 18340 12292
rect 18060 11788 18116 11844
rect 18956 14812 19012 14868
rect 18620 12962 18676 12964
rect 18620 12910 18622 12962
rect 18622 12910 18674 12962
rect 18674 12910 18676 12962
rect 18620 12908 18676 12910
rect 18508 12850 18564 12852
rect 18508 12798 18510 12850
rect 18510 12798 18562 12850
rect 18562 12798 18564 12850
rect 18508 12796 18564 12798
rect 18508 12402 18564 12404
rect 18508 12350 18510 12402
rect 18510 12350 18562 12402
rect 18562 12350 18564 12402
rect 18508 12348 18564 12350
rect 19516 16828 19572 16884
rect 20412 21586 20468 21588
rect 20412 21534 20414 21586
rect 20414 21534 20466 21586
rect 20466 21534 20468 21586
rect 20412 21532 20468 21534
rect 20636 23826 20692 23828
rect 20636 23774 20638 23826
rect 20638 23774 20690 23826
rect 20690 23774 20692 23826
rect 20636 23772 20692 23774
rect 22092 26348 22148 26404
rect 22652 26290 22708 26292
rect 22652 26238 22654 26290
rect 22654 26238 22706 26290
rect 22706 26238 22708 26290
rect 22652 26236 22708 26238
rect 21308 25394 21364 25396
rect 21308 25342 21310 25394
rect 21310 25342 21362 25394
rect 21362 25342 21364 25394
rect 21308 25340 21364 25342
rect 21196 24610 21252 24612
rect 21196 24558 21198 24610
rect 21198 24558 21250 24610
rect 21250 24558 21252 24610
rect 21196 24556 21252 24558
rect 21644 24556 21700 24612
rect 21980 24332 22036 24388
rect 22092 26012 22148 26068
rect 21868 24220 21924 24276
rect 22672 25898 22728 25900
rect 22672 25846 22674 25898
rect 22674 25846 22726 25898
rect 22726 25846 22728 25898
rect 22672 25844 22728 25846
rect 22776 25898 22832 25900
rect 22776 25846 22778 25898
rect 22778 25846 22830 25898
rect 22830 25846 22832 25898
rect 22776 25844 22832 25846
rect 22880 25898 22936 25900
rect 22880 25846 22882 25898
rect 22882 25846 22934 25898
rect 22934 25846 22936 25898
rect 22880 25844 22936 25846
rect 23100 25788 23156 25844
rect 22540 24722 22596 24724
rect 22540 24670 22542 24722
rect 22542 24670 22594 24722
rect 22594 24670 22596 24722
rect 22540 24668 22596 24670
rect 22204 24556 22260 24612
rect 22316 24220 22372 24276
rect 22428 24332 22484 24388
rect 22204 24108 22260 24164
rect 21868 23436 21924 23492
rect 21980 23772 22036 23828
rect 21420 23324 21476 23380
rect 21532 23212 21588 23268
rect 20860 22652 20916 22708
rect 20748 21756 20804 21812
rect 20860 22092 20916 22148
rect 21532 21756 21588 21812
rect 21420 21644 21476 21700
rect 20636 21420 20692 21476
rect 20748 20802 20804 20804
rect 20748 20750 20750 20802
rect 20750 20750 20802 20802
rect 20802 20750 20804 20802
rect 20748 20748 20804 20750
rect 20524 20188 20580 20244
rect 21420 20636 21476 20692
rect 21308 20018 21364 20020
rect 21308 19966 21310 20018
rect 21310 19966 21362 20018
rect 21362 19966 21364 20018
rect 21308 19964 21364 19966
rect 20412 17836 20468 17892
rect 20524 19852 20580 19908
rect 19740 16770 19796 16772
rect 19740 16718 19742 16770
rect 19742 16718 19794 16770
rect 19794 16718 19796 16770
rect 19740 16716 19796 16718
rect 20076 16098 20132 16100
rect 20076 16046 20078 16098
rect 20078 16046 20130 16098
rect 20130 16046 20132 16098
rect 20076 16044 20132 16046
rect 19404 14588 19460 14644
rect 19628 14476 19684 14532
rect 19068 13916 19124 13972
rect 21084 19516 21140 19572
rect 21532 20412 21588 20468
rect 20636 18844 20692 18900
rect 20748 18450 20804 18452
rect 20748 18398 20750 18450
rect 20750 18398 20802 18450
rect 20802 18398 20804 18450
rect 20748 18396 20804 18398
rect 21308 18396 21364 18452
rect 20412 16882 20468 16884
rect 20412 16830 20414 16882
rect 20414 16830 20466 16882
rect 20466 16830 20468 16882
rect 20412 16828 20468 16830
rect 20748 16492 20804 16548
rect 20300 14812 20356 14868
rect 20412 16268 20468 16324
rect 19292 13074 19348 13076
rect 19292 13022 19294 13074
rect 19294 13022 19346 13074
rect 19346 13022 19348 13074
rect 19292 13020 19348 13022
rect 19740 13020 19796 13076
rect 20636 13074 20692 13076
rect 20636 13022 20638 13074
rect 20638 13022 20690 13074
rect 20690 13022 20692 13074
rect 20636 13020 20692 13022
rect 20188 12962 20244 12964
rect 20188 12910 20190 12962
rect 20190 12910 20242 12962
rect 20242 12910 20244 12962
rect 20188 12908 20244 12910
rect 19964 12684 20020 12740
rect 18844 12402 18900 12404
rect 18844 12350 18846 12402
rect 18846 12350 18898 12402
rect 18898 12350 18900 12402
rect 18844 12348 18900 12350
rect 19180 12178 19236 12180
rect 19180 12126 19182 12178
rect 19182 12126 19234 12178
rect 19234 12126 19236 12178
rect 19180 12124 19236 12126
rect 18844 11788 18900 11844
rect 18284 10668 18340 10724
rect 19292 10722 19348 10724
rect 19292 10670 19294 10722
rect 19294 10670 19346 10722
rect 19346 10670 19348 10722
rect 19292 10668 19348 10670
rect 17612 10610 17668 10612
rect 17612 10558 17614 10610
rect 17614 10558 17666 10610
rect 17666 10558 17668 10610
rect 17612 10556 17668 10558
rect 17052 10444 17108 10500
rect 16268 9548 16324 9604
rect 17836 10386 17892 10388
rect 17836 10334 17838 10386
rect 17838 10334 17890 10386
rect 17890 10334 17892 10386
rect 17836 10332 17892 10334
rect 16828 9772 16884 9828
rect 18060 9772 18116 9828
rect 18284 9938 18340 9940
rect 18284 9886 18286 9938
rect 18286 9886 18338 9938
rect 18338 9886 18340 9938
rect 18284 9884 18340 9886
rect 17836 9714 17892 9716
rect 17836 9662 17838 9714
rect 17838 9662 17890 9714
rect 17890 9662 17892 9714
rect 17836 9660 17892 9662
rect 18956 9884 19012 9940
rect 19180 9772 19236 9828
rect 18844 9714 18900 9716
rect 18844 9662 18846 9714
rect 18846 9662 18898 9714
rect 18898 9662 18900 9714
rect 18844 9660 18900 9662
rect 17724 9154 17780 9156
rect 17724 9102 17726 9154
rect 17726 9102 17778 9154
rect 17778 9102 17780 9154
rect 17724 9100 17780 9102
rect 16716 8876 16772 8932
rect 17836 8876 17892 8932
rect 15932 8540 15988 8596
rect 16380 8540 16436 8596
rect 15596 8204 15652 8260
rect 15708 8146 15764 8148
rect 15708 8094 15710 8146
rect 15710 8094 15762 8146
rect 15762 8094 15764 8146
rect 15708 8092 15764 8094
rect 15518 7866 15574 7868
rect 15518 7814 15520 7866
rect 15520 7814 15572 7866
rect 15572 7814 15574 7866
rect 15518 7812 15574 7814
rect 15622 7866 15678 7868
rect 15622 7814 15624 7866
rect 15624 7814 15676 7866
rect 15676 7814 15678 7866
rect 15622 7812 15678 7814
rect 15726 7866 15782 7868
rect 15726 7814 15728 7866
rect 15728 7814 15780 7866
rect 15780 7814 15782 7866
rect 15726 7812 15782 7814
rect 15932 7084 15988 7140
rect 16044 6748 16100 6804
rect 15518 6298 15574 6300
rect 15518 6246 15520 6298
rect 15520 6246 15572 6298
rect 15572 6246 15574 6298
rect 15518 6244 15574 6246
rect 15622 6298 15678 6300
rect 15622 6246 15624 6298
rect 15624 6246 15676 6298
rect 15676 6246 15678 6298
rect 15622 6244 15678 6246
rect 15726 6298 15782 6300
rect 15726 6246 15728 6298
rect 15728 6246 15780 6298
rect 15780 6246 15782 6298
rect 15726 6244 15782 6246
rect 14812 5964 14868 6020
rect 15596 5404 15652 5460
rect 12908 4956 12964 5012
rect 12796 4508 12852 4564
rect 11788 4396 11844 4452
rect 13468 4562 13524 4564
rect 13468 4510 13470 4562
rect 13470 4510 13522 4562
rect 13522 4510 13524 4562
rect 13468 4508 13524 4510
rect 12012 4338 12068 4340
rect 12012 4286 12014 4338
rect 12014 4286 12066 4338
rect 12066 4286 12068 4338
rect 12012 4284 12068 4286
rect 12460 4338 12516 4340
rect 12460 4286 12462 4338
rect 12462 4286 12514 4338
rect 12514 4286 12516 4338
rect 12460 4284 12516 4286
rect 11452 4226 11508 4228
rect 11452 4174 11454 4226
rect 11454 4174 11506 4226
rect 11506 4174 11508 4226
rect 11452 4172 11508 4174
rect 13132 4172 13188 4228
rect 8365 3946 8421 3948
rect 8365 3894 8367 3946
rect 8367 3894 8419 3946
rect 8419 3894 8421 3946
rect 8365 3892 8421 3894
rect 8469 3946 8525 3948
rect 8469 3894 8471 3946
rect 8471 3894 8523 3946
rect 8523 3894 8525 3946
rect 8469 3892 8525 3894
rect 8573 3946 8629 3948
rect 8573 3894 8575 3946
rect 8575 3894 8627 3946
rect 8627 3894 8629 3946
rect 8573 3892 8629 3894
rect 13356 4338 13412 4340
rect 13356 4286 13358 4338
rect 13358 4286 13410 4338
rect 13410 4286 13412 4338
rect 13356 4284 13412 4286
rect 13804 5068 13860 5124
rect 18284 8428 18340 8484
rect 17500 6802 17556 6804
rect 17500 6750 17502 6802
rect 17502 6750 17554 6802
rect 17554 6750 17556 6802
rect 17500 6748 17556 6750
rect 18172 6748 18228 6804
rect 17388 6690 17444 6692
rect 17388 6638 17390 6690
rect 17390 6638 17442 6690
rect 17442 6638 17444 6690
rect 17388 6636 17444 6638
rect 18284 6636 18340 6692
rect 18508 7474 18564 7476
rect 18508 7422 18510 7474
rect 18510 7422 18562 7474
rect 18562 7422 18564 7474
rect 18508 7420 18564 7422
rect 21532 17612 21588 17668
rect 21420 17500 21476 17556
rect 20972 15932 21028 15988
rect 21084 16156 21140 16212
rect 22204 23826 22260 23828
rect 22204 23774 22206 23826
rect 22206 23774 22258 23826
rect 22258 23774 22260 23826
rect 22204 23772 22260 23774
rect 22652 24444 22708 24500
rect 22672 24330 22728 24332
rect 22672 24278 22674 24330
rect 22674 24278 22726 24330
rect 22726 24278 22728 24330
rect 22672 24276 22728 24278
rect 22776 24330 22832 24332
rect 22776 24278 22778 24330
rect 22778 24278 22830 24330
rect 22830 24278 22832 24330
rect 22776 24276 22832 24278
rect 22880 24330 22936 24332
rect 22880 24278 22882 24330
rect 22882 24278 22934 24330
rect 22934 24278 22936 24330
rect 22880 24276 22936 24278
rect 22540 23772 22596 23828
rect 22764 24108 22820 24164
rect 22428 23660 22484 23716
rect 22540 23548 22596 23604
rect 21868 22540 21924 22596
rect 22316 23378 22372 23380
rect 22316 23326 22318 23378
rect 22318 23326 22370 23378
rect 22370 23326 22372 23378
rect 22316 23324 22372 23326
rect 24668 26178 24724 26180
rect 24668 26126 24670 26178
rect 24670 26126 24722 26178
rect 24722 26126 24724 26178
rect 24668 26124 24724 26126
rect 23660 26066 23716 26068
rect 23660 26014 23662 26066
rect 23662 26014 23714 26066
rect 23714 26014 23716 26066
rect 23660 26012 23716 26014
rect 23996 26066 24052 26068
rect 23996 26014 23998 26066
rect 23998 26014 24050 26066
rect 24050 26014 24052 26066
rect 23996 26012 24052 26014
rect 25452 26178 25508 26180
rect 25452 26126 25454 26178
rect 25454 26126 25506 26178
rect 25506 26126 25508 26178
rect 25452 26124 25508 26126
rect 25228 26012 25284 26068
rect 26012 25788 26068 25844
rect 26236 25788 26292 25844
rect 23436 24780 23492 24836
rect 24668 24834 24724 24836
rect 24668 24782 24670 24834
rect 24670 24782 24722 24834
rect 24722 24782 24724 24834
rect 24668 24780 24724 24782
rect 24444 24444 24500 24500
rect 24780 23772 24836 23828
rect 23324 23436 23380 23492
rect 22204 22316 22260 22372
rect 22672 22762 22728 22764
rect 22672 22710 22674 22762
rect 22674 22710 22726 22762
rect 22726 22710 22728 22762
rect 22672 22708 22728 22710
rect 22776 22762 22832 22764
rect 22776 22710 22778 22762
rect 22778 22710 22830 22762
rect 22830 22710 22832 22762
rect 22776 22708 22832 22710
rect 22880 22762 22936 22764
rect 22880 22710 22882 22762
rect 22882 22710 22934 22762
rect 22934 22710 22936 22762
rect 22880 22708 22936 22710
rect 22988 22540 23044 22596
rect 22540 22204 22596 22260
rect 22204 21532 22260 21588
rect 22428 21980 22484 22036
rect 22764 22146 22820 22148
rect 22764 22094 22766 22146
rect 22766 22094 22818 22146
rect 22818 22094 22820 22146
rect 22764 22092 22820 22094
rect 23884 23154 23940 23156
rect 23884 23102 23886 23154
rect 23886 23102 23938 23154
rect 23938 23102 23940 23154
rect 23884 23100 23940 23102
rect 22672 21194 22728 21196
rect 22672 21142 22674 21194
rect 22674 21142 22726 21194
rect 22726 21142 22728 21194
rect 22672 21140 22728 21142
rect 22776 21194 22832 21196
rect 22776 21142 22778 21194
rect 22778 21142 22830 21194
rect 22830 21142 22832 21194
rect 22776 21140 22832 21142
rect 22880 21194 22936 21196
rect 22880 21142 22882 21194
rect 22882 21142 22934 21194
rect 22934 21142 22936 21194
rect 22880 21140 22936 21142
rect 22540 20748 22596 20804
rect 23324 20802 23380 20804
rect 23324 20750 23326 20802
rect 23326 20750 23378 20802
rect 23378 20750 23380 20802
rect 23324 20748 23380 20750
rect 22652 20578 22708 20580
rect 22652 20526 22654 20578
rect 22654 20526 22706 20578
rect 22706 20526 22708 20578
rect 22652 20524 22708 20526
rect 23548 22316 23604 22372
rect 23884 21586 23940 21588
rect 23884 21534 23886 21586
rect 23886 21534 23938 21586
rect 23938 21534 23940 21586
rect 23884 21532 23940 21534
rect 24444 23436 24500 23492
rect 25340 24444 25396 24500
rect 24556 23378 24612 23380
rect 24556 23326 24558 23378
rect 24558 23326 24610 23378
rect 24610 23326 24612 23378
rect 24556 23324 24612 23326
rect 24668 22594 24724 22596
rect 24668 22542 24670 22594
rect 24670 22542 24722 22594
rect 24722 22542 24724 22594
rect 24668 22540 24724 22542
rect 24332 22204 24388 22260
rect 23996 21196 24052 21252
rect 24556 21196 24612 21252
rect 21868 19852 21924 19908
rect 22672 19626 22728 19628
rect 22672 19574 22674 19626
rect 22674 19574 22726 19626
rect 22726 19574 22728 19626
rect 22672 19572 22728 19574
rect 22776 19626 22832 19628
rect 22776 19574 22778 19626
rect 22778 19574 22830 19626
rect 22830 19574 22832 19626
rect 22776 19572 22832 19574
rect 22880 19626 22936 19628
rect 22880 19574 22882 19626
rect 22882 19574 22934 19626
rect 22934 19574 22936 19626
rect 22880 19572 22936 19574
rect 23548 19516 23604 19572
rect 22204 18956 22260 19012
rect 22092 18508 22148 18564
rect 21868 17836 21924 17892
rect 21532 16044 21588 16100
rect 21980 15986 22036 15988
rect 21980 15934 21982 15986
rect 21982 15934 22034 15986
rect 22034 15934 22036 15986
rect 21980 15932 22036 15934
rect 21196 13804 21252 13860
rect 21084 13692 21140 13748
rect 20748 11394 20804 11396
rect 20748 11342 20750 11394
rect 20750 11342 20802 11394
rect 20802 11342 20804 11394
rect 20748 11340 20804 11342
rect 22540 18508 22596 18564
rect 22764 18284 22820 18340
rect 22672 18058 22728 18060
rect 22672 18006 22674 18058
rect 22674 18006 22726 18058
rect 22726 18006 22728 18058
rect 22672 18004 22728 18006
rect 22776 18058 22832 18060
rect 22776 18006 22778 18058
rect 22778 18006 22830 18058
rect 22830 18006 22832 18058
rect 22776 18004 22832 18006
rect 22880 18058 22936 18060
rect 22880 18006 22882 18058
rect 22882 18006 22934 18058
rect 22934 18006 22936 18058
rect 22880 18004 22936 18006
rect 23100 17836 23156 17892
rect 23212 18956 23268 19012
rect 23436 18508 23492 18564
rect 23212 17500 23268 17556
rect 23324 18284 23380 18340
rect 22428 16940 22484 16996
rect 22204 16098 22260 16100
rect 22204 16046 22206 16098
rect 22206 16046 22258 16098
rect 22258 16046 22260 16098
rect 22204 16044 22260 16046
rect 23324 16994 23380 16996
rect 23324 16942 23326 16994
rect 23326 16942 23378 16994
rect 23378 16942 23380 16994
rect 23324 16940 23380 16942
rect 23212 16716 23268 16772
rect 22672 16490 22728 16492
rect 22672 16438 22674 16490
rect 22674 16438 22726 16490
rect 22726 16438 22728 16490
rect 22672 16436 22728 16438
rect 22776 16490 22832 16492
rect 22776 16438 22778 16490
rect 22778 16438 22830 16490
rect 22830 16438 22832 16490
rect 22776 16436 22832 16438
rect 22880 16490 22936 16492
rect 22880 16438 22882 16490
rect 22882 16438 22934 16490
rect 22934 16438 22936 16490
rect 22880 16436 22936 16438
rect 22316 15820 22372 15876
rect 22428 15148 22484 15204
rect 21532 14588 21588 14644
rect 21868 14476 21924 14532
rect 23212 16098 23268 16100
rect 23212 16046 23214 16098
rect 23214 16046 23266 16098
rect 23266 16046 23268 16098
rect 23212 16044 23268 16046
rect 23548 17164 23604 17220
rect 23436 16156 23492 16212
rect 22672 14922 22728 14924
rect 22672 14870 22674 14922
rect 22674 14870 22726 14922
rect 22726 14870 22728 14922
rect 22672 14868 22728 14870
rect 22776 14922 22832 14924
rect 22776 14870 22778 14922
rect 22778 14870 22830 14922
rect 22830 14870 22832 14922
rect 22776 14868 22832 14870
rect 22880 14922 22936 14924
rect 22880 14870 22882 14922
rect 22882 14870 22934 14922
rect 22934 14870 22936 14922
rect 22880 14868 22936 14870
rect 23324 14476 23380 14532
rect 23436 14924 23492 14980
rect 22988 14140 23044 14196
rect 21644 13804 21700 13860
rect 22204 13522 22260 13524
rect 22204 13470 22206 13522
rect 22206 13470 22258 13522
rect 22258 13470 22260 13522
rect 22204 13468 22260 13470
rect 23100 13804 23156 13860
rect 23772 19516 23828 19572
rect 24668 19964 24724 20020
rect 24556 19404 24612 19460
rect 24220 18396 24276 18452
rect 24668 18338 24724 18340
rect 24668 18286 24670 18338
rect 24670 18286 24722 18338
rect 24722 18286 24724 18338
rect 24668 18284 24724 18286
rect 24332 17554 24388 17556
rect 24332 17502 24334 17554
rect 24334 17502 24386 17554
rect 24386 17502 24388 17554
rect 24332 17500 24388 17502
rect 23772 17052 23828 17108
rect 24444 17052 24500 17108
rect 24332 16658 24388 16660
rect 24332 16606 24334 16658
rect 24334 16606 24386 16658
rect 24386 16606 24388 16658
rect 24332 16604 24388 16606
rect 23884 16044 23940 16100
rect 25228 22652 25284 22708
rect 25340 20748 25396 20804
rect 25228 19516 25284 19572
rect 25340 20524 25396 20580
rect 25004 18620 25060 18676
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 26460 25564 26516 25620
rect 25676 23324 25732 23380
rect 25788 23548 25844 23604
rect 25676 23042 25732 23044
rect 25676 22990 25678 23042
rect 25678 22990 25730 23042
rect 25730 22990 25732 23042
rect 25676 22988 25732 22990
rect 25676 21980 25732 22036
rect 28924 26402 28980 26404
rect 28924 26350 28926 26402
rect 28926 26350 28978 26402
rect 28978 26350 28980 26402
rect 28924 26348 28980 26350
rect 26236 23996 26292 24052
rect 27356 26290 27412 26292
rect 27356 26238 27358 26290
rect 27358 26238 27410 26290
rect 27410 26238 27412 26290
rect 27356 26236 27412 26238
rect 27020 25900 27076 25956
rect 26684 23660 26740 23716
rect 26348 23436 26404 23492
rect 26460 23042 26516 23044
rect 26460 22990 26462 23042
rect 26462 22990 26514 23042
rect 26514 22990 26516 23042
rect 26460 22988 26516 22990
rect 26796 22652 26852 22708
rect 26796 22258 26852 22260
rect 26796 22206 26798 22258
rect 26798 22206 26850 22258
rect 26850 22206 26852 22258
rect 26796 22204 26852 22206
rect 26572 21810 26628 21812
rect 26572 21758 26574 21810
rect 26574 21758 26626 21810
rect 26626 21758 26628 21810
rect 26572 21756 26628 21758
rect 26124 21644 26180 21700
rect 25676 21474 25732 21476
rect 25676 21422 25678 21474
rect 25678 21422 25730 21474
rect 25730 21422 25732 21474
rect 25676 21420 25732 21422
rect 28700 26290 28756 26292
rect 28700 26238 28702 26290
rect 28702 26238 28754 26290
rect 28754 26238 28756 26290
rect 28700 26236 28756 26238
rect 27356 25788 27412 25844
rect 28476 25394 28532 25396
rect 28476 25342 28478 25394
rect 28478 25342 28530 25394
rect 28530 25342 28532 25394
rect 28476 25340 28532 25342
rect 27132 23436 27188 23492
rect 27020 23324 27076 23380
rect 28364 24722 28420 24724
rect 28364 24670 28366 24722
rect 28366 24670 28418 24722
rect 28418 24670 28420 24722
rect 28364 24668 28420 24670
rect 27804 23938 27860 23940
rect 27804 23886 27806 23938
rect 27806 23886 27858 23938
rect 27858 23886 27860 23938
rect 27804 23884 27860 23886
rect 27020 21532 27076 21588
rect 26348 20188 26404 20244
rect 25900 20018 25956 20020
rect 25900 19966 25902 20018
rect 25902 19966 25954 20018
rect 25954 19966 25956 20018
rect 25900 19964 25956 19966
rect 26236 19458 26292 19460
rect 26236 19406 26238 19458
rect 26238 19406 26290 19458
rect 26290 19406 26292 19458
rect 26236 19404 26292 19406
rect 26124 19292 26180 19348
rect 25900 18956 25956 19012
rect 25900 18620 25956 18676
rect 25340 17948 25396 18004
rect 25564 18284 25620 18340
rect 25340 17442 25396 17444
rect 25340 17390 25342 17442
rect 25342 17390 25394 17442
rect 25394 17390 25396 17442
rect 25340 17388 25396 17390
rect 26236 19068 26292 19124
rect 26572 20076 26628 20132
rect 27020 19068 27076 19124
rect 26460 18956 26516 19012
rect 26908 18844 26964 18900
rect 26572 18508 26628 18564
rect 25564 16940 25620 16996
rect 24780 16492 24836 16548
rect 24556 16098 24612 16100
rect 24556 16046 24558 16098
rect 24558 16046 24610 16098
rect 24610 16046 24612 16098
rect 24556 16044 24612 16046
rect 25452 16044 25508 16100
rect 24556 15820 24612 15876
rect 24108 15202 24164 15204
rect 24108 15150 24110 15202
rect 24110 15150 24162 15202
rect 24162 15150 24164 15202
rect 24108 15148 24164 15150
rect 26460 17724 26516 17780
rect 26012 17500 26068 17556
rect 26236 17388 26292 17444
rect 26460 17052 26516 17108
rect 26348 16882 26404 16884
rect 26348 16830 26350 16882
rect 26350 16830 26402 16882
rect 26402 16830 26404 16882
rect 26348 16828 26404 16830
rect 26124 16380 26180 16436
rect 27692 21586 27748 21588
rect 27692 21534 27694 21586
rect 27694 21534 27746 21586
rect 27746 21534 27748 21586
rect 27692 21532 27748 21534
rect 27468 19292 27524 19348
rect 27692 18844 27748 18900
rect 27356 18450 27412 18452
rect 27356 18398 27358 18450
rect 27358 18398 27410 18450
rect 27410 18398 27412 18450
rect 27356 18396 27412 18398
rect 28028 22652 28084 22708
rect 28252 20636 28308 20692
rect 28588 23884 28644 23940
rect 28700 23660 28756 23716
rect 28588 22652 28644 22708
rect 29372 25618 29428 25620
rect 29372 25566 29374 25618
rect 29374 25566 29426 25618
rect 29426 25566 29428 25618
rect 29372 25564 29428 25566
rect 29825 26682 29881 26684
rect 29825 26630 29827 26682
rect 29827 26630 29879 26682
rect 29879 26630 29881 26682
rect 29825 26628 29881 26630
rect 29929 26682 29985 26684
rect 29929 26630 29931 26682
rect 29931 26630 29983 26682
rect 29983 26630 29985 26682
rect 29929 26628 29985 26630
rect 30033 26682 30089 26684
rect 30033 26630 30035 26682
rect 30035 26630 30087 26682
rect 30087 26630 30089 26682
rect 30033 26628 30089 26630
rect 44132 26682 44188 26684
rect 44132 26630 44134 26682
rect 44134 26630 44186 26682
rect 44186 26630 44188 26682
rect 44132 26628 44188 26630
rect 44236 26682 44292 26684
rect 44236 26630 44238 26682
rect 44238 26630 44290 26682
rect 44290 26630 44292 26682
rect 44236 26628 44292 26630
rect 44340 26682 44396 26684
rect 44340 26630 44342 26682
rect 44342 26630 44394 26682
rect 44394 26630 44396 26682
rect 44340 26628 44396 26630
rect 29932 26348 29988 26404
rect 36092 26348 36148 26404
rect 29820 25564 29876 25620
rect 31276 26290 31332 26292
rect 31276 26238 31278 26290
rect 31278 26238 31330 26290
rect 31330 26238 31332 26290
rect 31276 26236 31332 26238
rect 29825 25114 29881 25116
rect 29825 25062 29827 25114
rect 29827 25062 29879 25114
rect 29879 25062 29881 25114
rect 29825 25060 29881 25062
rect 29929 25114 29985 25116
rect 29929 25062 29931 25114
rect 29931 25062 29983 25114
rect 29983 25062 29985 25114
rect 29929 25060 29985 25062
rect 30033 25114 30089 25116
rect 30033 25062 30035 25114
rect 30035 25062 30087 25114
rect 30087 25062 30089 25114
rect 30033 25060 30089 25062
rect 29596 24892 29652 24948
rect 29596 24668 29652 24724
rect 29260 23826 29316 23828
rect 29260 23774 29262 23826
rect 29262 23774 29314 23826
rect 29314 23774 29316 23826
rect 29260 23772 29316 23774
rect 29148 23548 29204 23604
rect 28924 22876 28980 22932
rect 30604 24892 30660 24948
rect 29825 23546 29881 23548
rect 29825 23494 29827 23546
rect 29827 23494 29879 23546
rect 29879 23494 29881 23546
rect 29825 23492 29881 23494
rect 29929 23546 29985 23548
rect 29929 23494 29931 23546
rect 29931 23494 29983 23546
rect 29983 23494 29985 23546
rect 29929 23492 29985 23494
rect 30033 23546 30089 23548
rect 30033 23494 30035 23546
rect 30035 23494 30087 23546
rect 30087 23494 30089 23546
rect 30033 23492 30089 23494
rect 29708 23100 29764 23156
rect 30492 24722 30548 24724
rect 30492 24670 30494 24722
rect 30494 24670 30546 24722
rect 30546 24670 30548 24722
rect 30492 24668 30548 24670
rect 31164 25116 31220 25172
rect 31052 24780 31108 24836
rect 31948 25900 32004 25956
rect 31612 25564 31668 25620
rect 31388 24946 31444 24948
rect 31388 24894 31390 24946
rect 31390 24894 31442 24946
rect 31442 24894 31444 24946
rect 31388 24892 31444 24894
rect 31388 24668 31444 24724
rect 30380 23436 30436 23492
rect 31052 23324 31108 23380
rect 30492 23042 30548 23044
rect 30492 22990 30494 23042
rect 30494 22990 30546 23042
rect 30546 22990 30548 23042
rect 30492 22988 30548 22990
rect 30380 22876 30436 22932
rect 29825 21978 29881 21980
rect 29825 21926 29827 21978
rect 29827 21926 29879 21978
rect 29879 21926 29881 21978
rect 29825 21924 29881 21926
rect 29929 21978 29985 21980
rect 29929 21926 29931 21978
rect 29931 21926 29983 21978
rect 29983 21926 29985 21978
rect 29929 21924 29985 21926
rect 30033 21978 30089 21980
rect 30033 21926 30035 21978
rect 30035 21926 30087 21978
rect 30087 21926 30089 21978
rect 30033 21924 30089 21926
rect 30380 21756 30436 21812
rect 28476 21420 28532 21476
rect 27916 18284 27972 18340
rect 29148 20188 29204 20244
rect 28476 19180 28532 19236
rect 28028 17836 28084 17892
rect 29372 20690 29428 20692
rect 29372 20638 29374 20690
rect 29374 20638 29426 20690
rect 29426 20638 29428 20690
rect 29372 20636 29428 20638
rect 29820 20690 29876 20692
rect 29820 20638 29822 20690
rect 29822 20638 29874 20690
rect 29874 20638 29876 20690
rect 29820 20636 29876 20638
rect 29825 20410 29881 20412
rect 29825 20358 29827 20410
rect 29827 20358 29879 20410
rect 29879 20358 29881 20410
rect 29825 20356 29881 20358
rect 29929 20410 29985 20412
rect 29929 20358 29931 20410
rect 29931 20358 29983 20410
rect 29983 20358 29985 20410
rect 29929 20356 29985 20358
rect 30033 20410 30089 20412
rect 30033 20358 30035 20410
rect 30035 20358 30087 20410
rect 30087 20358 30089 20410
rect 30033 20356 30089 20358
rect 30156 20188 30212 20244
rect 30268 21196 30324 21252
rect 29484 19794 29540 19796
rect 29484 19742 29486 19794
rect 29486 19742 29538 19794
rect 29538 19742 29540 19794
rect 29484 19740 29540 19742
rect 28588 18620 28644 18676
rect 28700 18508 28756 18564
rect 30044 19292 30100 19348
rect 31388 22988 31444 23044
rect 30604 20636 30660 20692
rect 29825 18842 29881 18844
rect 29825 18790 29827 18842
rect 29827 18790 29879 18842
rect 29879 18790 29881 18842
rect 29825 18788 29881 18790
rect 29929 18842 29985 18844
rect 29929 18790 29931 18842
rect 29931 18790 29983 18842
rect 29983 18790 29985 18842
rect 29929 18788 29985 18790
rect 30033 18842 30089 18844
rect 30033 18790 30035 18842
rect 30035 18790 30087 18842
rect 30087 18790 30089 18842
rect 30033 18788 30089 18790
rect 29708 18508 29764 18564
rect 29148 18450 29204 18452
rect 29148 18398 29150 18450
rect 29150 18398 29202 18450
rect 29202 18398 29204 18450
rect 29148 18396 29204 18398
rect 28364 17666 28420 17668
rect 28364 17614 28366 17666
rect 28366 17614 28418 17666
rect 28418 17614 28420 17666
rect 28364 17612 28420 17614
rect 27692 17554 27748 17556
rect 27692 17502 27694 17554
rect 27694 17502 27746 17554
rect 27746 17502 27748 17554
rect 27692 17500 27748 17502
rect 27356 17276 27412 17332
rect 28364 17164 28420 17220
rect 27244 16940 27300 16996
rect 27692 16882 27748 16884
rect 27692 16830 27694 16882
rect 27694 16830 27746 16882
rect 27746 16830 27748 16882
rect 27692 16828 27748 16830
rect 27020 16380 27076 16436
rect 26012 15820 26068 15876
rect 26684 15874 26740 15876
rect 26684 15822 26686 15874
rect 26686 15822 26738 15874
rect 26738 15822 26740 15874
rect 26684 15820 26740 15822
rect 26908 15708 26964 15764
rect 27132 16098 27188 16100
rect 27132 16046 27134 16098
rect 27134 16046 27186 16098
rect 27186 16046 27188 16098
rect 27132 16044 27188 16046
rect 27020 15484 27076 15540
rect 27916 16492 27972 16548
rect 28252 16492 28308 16548
rect 28140 16044 28196 16100
rect 27692 15708 27748 15764
rect 28588 15932 28644 15988
rect 28476 15874 28532 15876
rect 28476 15822 28478 15874
rect 28478 15822 28530 15874
rect 28530 15822 28532 15874
rect 28476 15820 28532 15822
rect 28364 15708 28420 15764
rect 24780 14924 24836 14980
rect 23884 14642 23940 14644
rect 23884 14590 23886 14642
rect 23886 14590 23938 14642
rect 23938 14590 23940 14642
rect 23884 14588 23940 14590
rect 23548 14476 23604 14532
rect 24444 14530 24500 14532
rect 24444 14478 24446 14530
rect 24446 14478 24498 14530
rect 24498 14478 24500 14530
rect 24444 14476 24500 14478
rect 25116 14588 25172 14644
rect 23772 14140 23828 14196
rect 28252 15260 28308 15316
rect 24780 13916 24836 13972
rect 21420 13356 21476 13412
rect 22672 13354 22728 13356
rect 22672 13302 22674 13354
rect 22674 13302 22726 13354
rect 22726 13302 22728 13354
rect 22672 13300 22728 13302
rect 22776 13354 22832 13356
rect 22776 13302 22778 13354
rect 22778 13302 22830 13354
rect 22830 13302 22832 13354
rect 22776 13300 22832 13302
rect 22880 13354 22936 13356
rect 22880 13302 22882 13354
rect 22882 13302 22934 13354
rect 22934 13302 22936 13354
rect 22880 13300 22936 13302
rect 22092 13132 22148 13188
rect 21868 12962 21924 12964
rect 21868 12910 21870 12962
rect 21870 12910 21922 12962
rect 21922 12910 21924 12962
rect 21868 12908 21924 12910
rect 21644 12066 21700 12068
rect 21644 12014 21646 12066
rect 21646 12014 21698 12066
rect 21698 12014 21700 12066
rect 21644 12012 21700 12014
rect 22988 13132 23044 13188
rect 22540 13020 22596 13076
rect 21980 12012 22036 12068
rect 22204 11900 22260 11956
rect 23212 13468 23268 13524
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 24332 13468 24388 13524
rect 23772 13132 23828 13188
rect 23324 13020 23380 13076
rect 23100 12348 23156 12404
rect 23100 12124 23156 12180
rect 22672 11786 22728 11788
rect 22672 11734 22674 11786
rect 22674 11734 22726 11786
rect 22726 11734 22728 11786
rect 22672 11732 22728 11734
rect 22776 11786 22832 11788
rect 22776 11734 22778 11786
rect 22778 11734 22830 11786
rect 22830 11734 22832 11786
rect 22776 11732 22832 11734
rect 22880 11786 22936 11788
rect 22880 11734 22882 11786
rect 22882 11734 22934 11786
rect 22934 11734 22936 11786
rect 22880 11732 22936 11734
rect 19964 10668 20020 10724
rect 19964 10332 20020 10388
rect 20748 10332 20804 10388
rect 21084 9100 21140 9156
rect 19628 8876 19684 8932
rect 20412 8876 20468 8932
rect 20188 8204 20244 8260
rect 18620 6748 18676 6804
rect 19068 7420 19124 7476
rect 18508 6690 18564 6692
rect 18508 6638 18510 6690
rect 18510 6638 18562 6690
rect 18562 6638 18564 6690
rect 18508 6636 18564 6638
rect 20188 7474 20244 7476
rect 20188 7422 20190 7474
rect 20190 7422 20242 7474
rect 20242 7422 20244 7474
rect 20188 7420 20244 7422
rect 21308 8876 21364 8932
rect 20524 8146 20580 8148
rect 20524 8094 20526 8146
rect 20526 8094 20578 8146
rect 20578 8094 20580 8146
rect 20524 8092 20580 8094
rect 21084 7474 21140 7476
rect 21084 7422 21086 7474
rect 21086 7422 21138 7474
rect 21138 7422 21140 7474
rect 21084 7420 21140 7422
rect 22316 11394 22372 11396
rect 22316 11342 22318 11394
rect 22318 11342 22370 11394
rect 22370 11342 22372 11394
rect 22316 11340 22372 11342
rect 21644 10722 21700 10724
rect 21644 10670 21646 10722
rect 21646 10670 21698 10722
rect 21698 10670 21700 10722
rect 21644 10668 21700 10670
rect 22428 10668 22484 10724
rect 21868 10332 21924 10388
rect 23436 11900 23492 11956
rect 23100 11282 23156 11284
rect 23100 11230 23102 11282
rect 23102 11230 23154 11282
rect 23154 11230 23156 11282
rect 23100 11228 23156 11230
rect 22876 10332 22932 10388
rect 22672 10218 22728 10220
rect 22672 10166 22674 10218
rect 22674 10166 22726 10218
rect 22726 10166 22728 10218
rect 22672 10164 22728 10166
rect 22776 10218 22832 10220
rect 22776 10166 22778 10218
rect 22778 10166 22830 10218
rect 22830 10166 22832 10218
rect 22776 10164 22832 10166
rect 22880 10218 22936 10220
rect 22880 10166 22882 10218
rect 22882 10166 22934 10218
rect 22934 10166 22936 10218
rect 22880 10164 22936 10166
rect 25900 13970 25956 13972
rect 25900 13918 25902 13970
rect 25902 13918 25954 13970
rect 25954 13918 25956 13970
rect 25900 13916 25956 13918
rect 25340 13746 25396 13748
rect 25340 13694 25342 13746
rect 25342 13694 25394 13746
rect 25394 13694 25396 13746
rect 25340 13692 25396 13694
rect 25228 13132 25284 13188
rect 23996 12348 24052 12404
rect 24668 12402 24724 12404
rect 24668 12350 24670 12402
rect 24670 12350 24722 12402
rect 24722 12350 24724 12402
rect 24668 12348 24724 12350
rect 25564 12348 25620 12404
rect 23772 11004 23828 11060
rect 23324 9772 23380 9828
rect 21980 9042 22036 9044
rect 21980 8990 21982 9042
rect 21982 8990 22034 9042
rect 22034 8990 22036 9042
rect 21980 8988 22036 8990
rect 21532 8258 21588 8260
rect 21532 8206 21534 8258
rect 21534 8206 21586 8258
rect 21586 8206 21588 8258
rect 21532 8204 21588 8206
rect 21868 8258 21924 8260
rect 21868 8206 21870 8258
rect 21870 8206 21922 8258
rect 21922 8206 21924 8258
rect 21868 8204 21924 8206
rect 22540 9154 22596 9156
rect 22540 9102 22542 9154
rect 22542 9102 22594 9154
rect 22594 9102 22596 9154
rect 22540 9100 22596 9102
rect 22672 8650 22728 8652
rect 22672 8598 22674 8650
rect 22674 8598 22726 8650
rect 22726 8598 22728 8650
rect 22672 8596 22728 8598
rect 22776 8650 22832 8652
rect 22776 8598 22778 8650
rect 22778 8598 22830 8650
rect 22830 8598 22832 8650
rect 22776 8596 22832 8598
rect 22880 8650 22936 8652
rect 22880 8598 22882 8650
rect 22882 8598 22934 8650
rect 22934 8598 22936 8650
rect 22880 8596 22936 8598
rect 23436 8204 23492 8260
rect 23436 7868 23492 7924
rect 22672 7082 22728 7084
rect 22672 7030 22674 7082
rect 22674 7030 22726 7082
rect 22726 7030 22728 7082
rect 22672 7028 22728 7030
rect 22776 7082 22832 7084
rect 22776 7030 22778 7082
rect 22778 7030 22830 7082
rect 22830 7030 22832 7082
rect 22776 7028 22832 7030
rect 22880 7082 22936 7084
rect 22880 7030 22882 7082
rect 22882 7030 22934 7082
rect 22934 7030 22936 7082
rect 22880 7028 22936 7030
rect 20524 6748 20580 6804
rect 19068 6076 19124 6132
rect 18508 5852 18564 5908
rect 18844 5906 18900 5908
rect 18844 5854 18846 5906
rect 18846 5854 18898 5906
rect 18898 5854 18900 5906
rect 18844 5852 18900 5854
rect 16156 5292 16212 5348
rect 15820 5010 15876 5012
rect 15820 4958 15822 5010
rect 15822 4958 15874 5010
rect 15874 4958 15876 5010
rect 15820 4956 15876 4958
rect 15518 4730 15574 4732
rect 15518 4678 15520 4730
rect 15520 4678 15572 4730
rect 15572 4678 15574 4730
rect 15518 4676 15574 4678
rect 15622 4730 15678 4732
rect 15622 4678 15624 4730
rect 15624 4678 15676 4730
rect 15676 4678 15678 4730
rect 15622 4676 15678 4678
rect 15726 4730 15782 4732
rect 15726 4678 15728 4730
rect 15728 4678 15780 4730
rect 15780 4678 15782 4730
rect 15726 4676 15782 4678
rect 13916 4284 13972 4340
rect 17948 5404 18004 5460
rect 16380 5122 16436 5124
rect 16380 5070 16382 5122
rect 16382 5070 16434 5122
rect 16434 5070 16436 5122
rect 16380 5068 16436 5070
rect 16716 4620 16772 4676
rect 16380 4450 16436 4452
rect 16380 4398 16382 4450
rect 16382 4398 16434 4450
rect 16434 4398 16436 4450
rect 16380 4396 16436 4398
rect 14476 4284 14532 4340
rect 19180 5404 19236 5460
rect 18732 4956 18788 5012
rect 18060 4450 18116 4452
rect 18060 4398 18062 4450
rect 18062 4398 18114 4450
rect 18114 4398 18116 4450
rect 18060 4396 18116 4398
rect 19628 4956 19684 5012
rect 19740 5404 19796 5460
rect 23884 6860 23940 6916
rect 21420 6748 21476 6804
rect 23324 6412 23380 6468
rect 21308 5852 21364 5908
rect 20636 4844 20692 4900
rect 20076 4450 20132 4452
rect 20076 4398 20078 4450
rect 20078 4398 20130 4450
rect 20130 4398 20132 4450
rect 20076 4396 20132 4398
rect 21644 5906 21700 5908
rect 21644 5854 21646 5906
rect 21646 5854 21698 5906
rect 21698 5854 21700 5906
rect 21644 5852 21700 5854
rect 21868 4956 21924 5012
rect 20972 4114 21028 4116
rect 20972 4062 20974 4114
rect 20974 4062 21026 4114
rect 21026 4062 21028 4114
rect 20972 4060 21028 4062
rect 19068 3724 19124 3780
rect 4284 3442 4340 3444
rect 4284 3390 4286 3442
rect 4286 3390 4338 3442
rect 4338 3390 4340 3442
rect 4284 3388 4340 3390
rect 22428 5906 22484 5908
rect 22428 5854 22430 5906
rect 22430 5854 22482 5906
rect 22482 5854 22484 5906
rect 22428 5852 22484 5854
rect 22672 5514 22728 5516
rect 22672 5462 22674 5514
rect 22674 5462 22726 5514
rect 22726 5462 22728 5514
rect 22672 5460 22728 5462
rect 22776 5514 22832 5516
rect 22776 5462 22778 5514
rect 22778 5462 22830 5514
rect 22830 5462 22832 5514
rect 22776 5460 22832 5462
rect 22880 5514 22936 5516
rect 22880 5462 22882 5514
rect 22882 5462 22934 5514
rect 22934 5462 22936 5514
rect 22880 5460 22936 5462
rect 22540 5234 22596 5236
rect 22540 5182 22542 5234
rect 22542 5182 22594 5234
rect 22594 5182 22596 5234
rect 22540 5180 22596 5182
rect 25228 11228 25284 11284
rect 24668 10834 24724 10836
rect 24668 10782 24670 10834
rect 24670 10782 24722 10834
rect 24722 10782 24724 10834
rect 24668 10780 24724 10782
rect 24444 9772 24500 9828
rect 24556 9100 24612 9156
rect 26796 14700 26852 14756
rect 28476 14588 28532 14644
rect 27468 14530 27524 14532
rect 27468 14478 27470 14530
rect 27470 14478 27522 14530
rect 27522 14478 27524 14530
rect 27468 14476 27524 14478
rect 28252 14476 28308 14532
rect 26796 14140 26852 14196
rect 27132 13916 27188 13972
rect 26124 13692 26180 13748
rect 26684 13746 26740 13748
rect 26684 13694 26686 13746
rect 26686 13694 26738 13746
rect 26738 13694 26740 13746
rect 26684 13692 26740 13694
rect 26236 12348 26292 12404
rect 26460 13468 26516 13524
rect 26908 13580 26964 13636
rect 27692 13970 27748 13972
rect 27692 13918 27694 13970
rect 27694 13918 27746 13970
rect 27746 13918 27748 13970
rect 27692 13916 27748 13918
rect 27804 13746 27860 13748
rect 27804 13694 27806 13746
rect 27806 13694 27858 13746
rect 27858 13694 27860 13746
rect 27804 13692 27860 13694
rect 31052 21586 31108 21588
rect 31052 21534 31054 21586
rect 31054 21534 31106 21586
rect 31106 21534 31108 21586
rect 31052 21532 31108 21534
rect 31052 20578 31108 20580
rect 31052 20526 31054 20578
rect 31054 20526 31106 20578
rect 31106 20526 31108 20578
rect 31052 20524 31108 20526
rect 30828 20300 30884 20356
rect 30716 19964 30772 20020
rect 32060 25452 32116 25508
rect 31836 25116 31892 25172
rect 31724 25004 31780 25060
rect 31612 20748 31668 20804
rect 31164 19234 31220 19236
rect 31164 19182 31166 19234
rect 31166 19182 31218 19234
rect 31218 19182 31220 19234
rect 31164 19180 31220 19182
rect 30380 17612 30436 17668
rect 29825 17274 29881 17276
rect 29825 17222 29827 17274
rect 29827 17222 29879 17274
rect 29879 17222 29881 17274
rect 29825 17220 29881 17222
rect 29929 17274 29985 17276
rect 29929 17222 29931 17274
rect 29931 17222 29983 17274
rect 29983 17222 29985 17274
rect 29929 17220 29985 17222
rect 30033 17274 30089 17276
rect 30033 17222 30035 17274
rect 30035 17222 30087 17274
rect 30087 17222 30089 17274
rect 30033 17220 30089 17222
rect 29260 16940 29316 16996
rect 29596 16882 29652 16884
rect 29596 16830 29598 16882
rect 29598 16830 29650 16882
rect 29650 16830 29652 16882
rect 29596 16828 29652 16830
rect 29596 16380 29652 16436
rect 31164 17612 31220 17668
rect 30716 16716 30772 16772
rect 30268 16492 30324 16548
rect 29825 15706 29881 15708
rect 29825 15654 29827 15706
rect 29827 15654 29879 15706
rect 29879 15654 29881 15706
rect 29825 15652 29881 15654
rect 29929 15706 29985 15708
rect 29929 15654 29931 15706
rect 29931 15654 29983 15706
rect 29983 15654 29985 15706
rect 29929 15652 29985 15654
rect 30033 15706 30089 15708
rect 30033 15654 30035 15706
rect 30035 15654 30087 15706
rect 30087 15654 30089 15706
rect 30033 15652 30089 15654
rect 30268 15484 30324 15540
rect 29825 14138 29881 14140
rect 29825 14086 29827 14138
rect 29827 14086 29879 14138
rect 29879 14086 29881 14138
rect 29825 14084 29881 14086
rect 29929 14138 29985 14140
rect 29929 14086 29931 14138
rect 29931 14086 29983 14138
rect 29983 14086 29985 14138
rect 29929 14084 29985 14086
rect 30033 14138 30089 14140
rect 30033 14086 30035 14138
rect 30035 14086 30087 14138
rect 30087 14086 30089 14138
rect 30033 14084 30089 14086
rect 28588 13804 28644 13860
rect 27916 13580 27972 13636
rect 30044 13858 30100 13860
rect 30044 13806 30046 13858
rect 30046 13806 30098 13858
rect 30098 13806 30100 13858
rect 30044 13804 30100 13806
rect 30828 15314 30884 15316
rect 30828 15262 30830 15314
rect 30830 15262 30882 15314
rect 30882 15262 30884 15314
rect 30828 15260 30884 15262
rect 28700 13580 28756 13636
rect 29708 13634 29764 13636
rect 29708 13582 29710 13634
rect 29710 13582 29762 13634
rect 29762 13582 29764 13634
rect 29708 13580 29764 13582
rect 27244 13132 27300 13188
rect 26460 12348 26516 12404
rect 25788 11282 25844 11284
rect 25788 11230 25790 11282
rect 25790 11230 25842 11282
rect 25842 11230 25844 11282
rect 25788 11228 25844 11230
rect 26796 11228 26852 11284
rect 26572 11116 26628 11172
rect 25900 11004 25956 11060
rect 25452 10610 25508 10612
rect 25452 10558 25454 10610
rect 25454 10558 25506 10610
rect 25506 10558 25508 10610
rect 25452 10556 25508 10558
rect 26572 10610 26628 10612
rect 26572 10558 26574 10610
rect 26574 10558 26626 10610
rect 26626 10558 26628 10610
rect 26572 10556 26628 10558
rect 26796 10556 26852 10612
rect 26908 10444 26964 10500
rect 26348 10332 26404 10388
rect 28252 13186 28308 13188
rect 28252 13134 28254 13186
rect 28254 13134 28306 13186
rect 28306 13134 28308 13186
rect 28252 13132 28308 13134
rect 29148 13132 29204 13188
rect 27692 12348 27748 12404
rect 28252 12348 28308 12404
rect 31164 14530 31220 14532
rect 31164 14478 31166 14530
rect 31166 14478 31218 14530
rect 31218 14478 31220 14530
rect 31164 14476 31220 14478
rect 30940 13186 30996 13188
rect 30940 13134 30942 13186
rect 30942 13134 30994 13186
rect 30994 13134 30996 13186
rect 30940 13132 30996 13134
rect 30716 12908 30772 12964
rect 31052 12908 31108 12964
rect 32396 25564 32452 25620
rect 32732 25452 32788 25508
rect 32172 24834 32228 24836
rect 32172 24782 32174 24834
rect 32174 24782 32226 24834
rect 32226 24782 32228 24834
rect 32172 24780 32228 24782
rect 31948 23436 32004 23492
rect 31836 20802 31892 20804
rect 31836 20750 31838 20802
rect 31838 20750 31890 20802
rect 31890 20750 31892 20802
rect 31836 20748 31892 20750
rect 32396 24780 32452 24836
rect 32844 25340 32900 25396
rect 33180 24668 33236 24724
rect 33180 24108 33236 24164
rect 33404 24834 33460 24836
rect 33404 24782 33406 24834
rect 33406 24782 33458 24834
rect 33458 24782 33460 24834
rect 33404 24780 33460 24782
rect 35532 26236 35588 26292
rect 34188 26124 34244 26180
rect 33740 25116 33796 25172
rect 33516 24668 33572 24724
rect 33404 23660 33460 23716
rect 32396 21196 32452 21252
rect 32172 20802 32228 20804
rect 32172 20750 32174 20802
rect 32174 20750 32226 20802
rect 32226 20750 32228 20802
rect 32172 20748 32228 20750
rect 32060 19180 32116 19236
rect 31948 18508 32004 18564
rect 31500 16492 31556 16548
rect 32060 17052 32116 17108
rect 32172 16828 32228 16884
rect 31724 16770 31780 16772
rect 31724 16718 31726 16770
rect 31726 16718 31778 16770
rect 31778 16718 31780 16770
rect 31724 16716 31780 16718
rect 31724 15202 31780 15204
rect 31724 15150 31726 15202
rect 31726 15150 31778 15202
rect 31778 15150 31780 15202
rect 31724 15148 31780 15150
rect 30604 12796 30660 12852
rect 27916 12066 27972 12068
rect 27916 12014 27918 12066
rect 27918 12014 27970 12066
rect 27970 12014 27972 12066
rect 27916 12012 27972 12014
rect 25788 9154 25844 9156
rect 25788 9102 25790 9154
rect 25790 9102 25842 9154
rect 25842 9102 25844 9154
rect 25788 9100 25844 9102
rect 26684 9154 26740 9156
rect 26684 9102 26686 9154
rect 26686 9102 26738 9154
rect 26738 9102 26740 9154
rect 26684 9100 26740 9102
rect 25004 8258 25060 8260
rect 25004 8206 25006 8258
rect 25006 8206 25058 8258
rect 25058 8206 25060 8258
rect 25004 8204 25060 8206
rect 25452 9042 25508 9044
rect 25452 8990 25454 9042
rect 25454 8990 25506 9042
rect 25506 8990 25508 9042
rect 25452 8988 25508 8990
rect 25676 8876 25732 8932
rect 24556 7644 24612 7700
rect 24332 6860 24388 6916
rect 22092 4508 22148 4564
rect 22876 4844 22932 4900
rect 22764 4450 22820 4452
rect 22764 4398 22766 4450
rect 22766 4398 22818 4450
rect 22818 4398 22820 4450
rect 22764 4396 22820 4398
rect 22428 4338 22484 4340
rect 22428 4286 22430 4338
rect 22430 4286 22482 4338
rect 22482 4286 22484 4338
rect 22428 4284 22484 4286
rect 21868 3778 21924 3780
rect 21868 3726 21870 3778
rect 21870 3726 21922 3778
rect 21922 3726 21924 3778
rect 21868 3724 21924 3726
rect 23996 4562 24052 4564
rect 23996 4510 23998 4562
rect 23998 4510 24050 4562
rect 24050 4510 24052 4562
rect 23996 4508 24052 4510
rect 25004 6860 25060 6916
rect 24780 6466 24836 6468
rect 24780 6414 24782 6466
rect 24782 6414 24834 6466
rect 24834 6414 24836 6466
rect 24780 6412 24836 6414
rect 24556 4620 24612 4676
rect 23772 4338 23828 4340
rect 23772 4286 23774 4338
rect 23774 4286 23826 4338
rect 23826 4286 23828 4338
rect 23772 4284 23828 4286
rect 23436 4114 23492 4116
rect 23436 4062 23438 4114
rect 23438 4062 23490 4114
rect 23490 4062 23492 4114
rect 23436 4060 23492 4062
rect 23772 4114 23828 4116
rect 23772 4062 23774 4114
rect 23774 4062 23826 4114
rect 23826 4062 23828 4114
rect 23772 4060 23828 4062
rect 22672 3946 22728 3948
rect 22672 3894 22674 3946
rect 22674 3894 22726 3946
rect 22726 3894 22728 3946
rect 22672 3892 22728 3894
rect 22776 3946 22832 3948
rect 22776 3894 22778 3946
rect 22778 3894 22830 3946
rect 22830 3894 22832 3946
rect 22776 3892 22832 3894
rect 22880 3946 22936 3948
rect 22880 3894 22882 3946
rect 22882 3894 22934 3946
rect 22934 3894 22936 3946
rect 24108 3948 24164 4004
rect 22880 3892 22936 3894
rect 23660 3724 23716 3780
rect 21084 3500 21140 3556
rect 21644 3554 21700 3556
rect 21644 3502 21646 3554
rect 21646 3502 21698 3554
rect 21698 3502 21700 3554
rect 21644 3500 21700 3502
rect 25452 7980 25508 8036
rect 26124 8988 26180 9044
rect 25900 8204 25956 8260
rect 26124 8204 26180 8260
rect 25788 8092 25844 8148
rect 25900 7868 25956 7924
rect 26124 7980 26180 8036
rect 25788 7586 25844 7588
rect 25788 7534 25790 7586
rect 25790 7534 25842 7586
rect 25842 7534 25844 7586
rect 25788 7532 25844 7534
rect 26572 8930 26628 8932
rect 26572 8878 26574 8930
rect 26574 8878 26626 8930
rect 26626 8878 26628 8930
rect 26572 8876 26628 8878
rect 27132 10668 27188 10724
rect 27356 9996 27412 10052
rect 28364 12178 28420 12180
rect 28364 12126 28366 12178
rect 28366 12126 28418 12178
rect 28418 12126 28420 12178
rect 28364 12124 28420 12126
rect 29825 12570 29881 12572
rect 29825 12518 29827 12570
rect 29827 12518 29879 12570
rect 29879 12518 29881 12570
rect 29825 12516 29881 12518
rect 29929 12570 29985 12572
rect 29929 12518 29931 12570
rect 29931 12518 29983 12570
rect 29983 12518 29985 12570
rect 29929 12516 29985 12518
rect 30033 12570 30089 12572
rect 30033 12518 30035 12570
rect 30035 12518 30087 12570
rect 30087 12518 30089 12570
rect 30033 12516 30089 12518
rect 29260 12124 29316 12180
rect 29148 11676 29204 11732
rect 28476 10668 28532 10724
rect 28812 11116 28868 11172
rect 30156 11618 30212 11620
rect 30156 11566 30158 11618
rect 30158 11566 30210 11618
rect 30210 11566 30212 11618
rect 30156 11564 30212 11566
rect 30380 11452 30436 11508
rect 30044 11282 30100 11284
rect 30044 11230 30046 11282
rect 30046 11230 30098 11282
rect 30098 11230 30100 11282
rect 30044 11228 30100 11230
rect 29820 11170 29876 11172
rect 29820 11118 29822 11170
rect 29822 11118 29874 11170
rect 29874 11118 29876 11170
rect 29820 11116 29876 11118
rect 29825 11002 29881 11004
rect 29825 10950 29827 11002
rect 29827 10950 29879 11002
rect 29879 10950 29881 11002
rect 29825 10948 29881 10950
rect 29929 11002 29985 11004
rect 29929 10950 29931 11002
rect 29931 10950 29983 11002
rect 29983 10950 29985 11002
rect 29929 10948 29985 10950
rect 30033 11002 30089 11004
rect 30033 10950 30035 11002
rect 30035 10950 30087 11002
rect 30087 10950 30089 11002
rect 30033 10948 30089 10950
rect 29484 10780 29540 10836
rect 29932 10834 29988 10836
rect 29932 10782 29934 10834
rect 29934 10782 29986 10834
rect 29986 10782 29988 10834
rect 29932 10780 29988 10782
rect 28812 10556 28868 10612
rect 31388 12908 31444 12964
rect 30380 10780 30436 10836
rect 28364 9996 28420 10052
rect 27468 9212 27524 9268
rect 27356 9154 27412 9156
rect 27356 9102 27358 9154
rect 27358 9102 27410 9154
rect 27410 9102 27412 9154
rect 27356 9100 27412 9102
rect 26908 8428 26964 8484
rect 26460 8258 26516 8260
rect 26460 8206 26462 8258
rect 26462 8206 26514 8258
rect 26514 8206 26516 8258
rect 26460 8204 26516 8206
rect 26236 7868 26292 7924
rect 26012 6748 26068 6804
rect 25676 5628 25732 5684
rect 25228 4620 25284 4676
rect 24668 3500 24724 3556
rect 23772 3442 23828 3444
rect 23772 3390 23774 3442
rect 23774 3390 23826 3442
rect 23826 3390 23828 3442
rect 23772 3388 23828 3390
rect 25788 5180 25844 5236
rect 28028 9212 28084 9268
rect 27132 8258 27188 8260
rect 27132 8206 27134 8258
rect 27134 8206 27186 8258
rect 27186 8206 27188 8258
rect 27132 8204 27188 8206
rect 28364 8316 28420 8372
rect 30716 9996 30772 10052
rect 32060 15820 32116 15876
rect 35420 26178 35476 26180
rect 35420 26126 35422 26178
rect 35422 26126 35474 26178
rect 35474 26126 35476 26178
rect 35420 26124 35476 26126
rect 35532 25618 35588 25620
rect 35532 25566 35534 25618
rect 35534 25566 35586 25618
rect 35586 25566 35588 25618
rect 35532 25564 35588 25566
rect 35980 26124 36036 26180
rect 34188 24780 34244 24836
rect 33740 23154 33796 23156
rect 33740 23102 33742 23154
rect 33742 23102 33794 23154
rect 33794 23102 33796 23154
rect 33740 23100 33796 23102
rect 33628 23042 33684 23044
rect 33628 22990 33630 23042
rect 33630 22990 33682 23042
rect 33682 22990 33684 23042
rect 33628 22988 33684 22990
rect 35420 25340 35476 25396
rect 34972 25282 35028 25284
rect 34972 25230 34974 25282
rect 34974 25230 35026 25282
rect 35026 25230 35028 25282
rect 34972 25228 35028 25230
rect 34972 24892 35028 24948
rect 34748 24780 34804 24836
rect 34524 24108 34580 24164
rect 34412 23100 34468 23156
rect 34748 24050 34804 24052
rect 34748 23998 34750 24050
rect 34750 23998 34802 24050
rect 34802 23998 34804 24050
rect 34748 23996 34804 23998
rect 35756 25116 35812 25172
rect 35420 23996 35476 24052
rect 35084 22876 35140 22932
rect 34412 21756 34468 21812
rect 35308 23714 35364 23716
rect 35308 23662 35310 23714
rect 35310 23662 35362 23714
rect 35362 23662 35364 23714
rect 35308 23660 35364 23662
rect 35308 23100 35364 23156
rect 36204 26290 36260 26292
rect 36204 26238 36206 26290
rect 36206 26238 36258 26290
rect 36258 26238 36260 26290
rect 36204 26236 36260 26238
rect 39116 26348 39172 26404
rect 37436 26012 37492 26068
rect 36979 25898 37035 25900
rect 36979 25846 36981 25898
rect 36981 25846 37033 25898
rect 37033 25846 37035 25898
rect 36979 25844 37035 25846
rect 37083 25898 37139 25900
rect 37083 25846 37085 25898
rect 37085 25846 37137 25898
rect 37137 25846 37139 25898
rect 37083 25844 37139 25846
rect 37187 25898 37243 25900
rect 37187 25846 37189 25898
rect 37189 25846 37241 25898
rect 37241 25846 37243 25898
rect 37187 25844 37243 25846
rect 36204 25452 36260 25508
rect 36428 25506 36484 25508
rect 36428 25454 36430 25506
rect 36430 25454 36482 25506
rect 36482 25454 36484 25506
rect 36428 25452 36484 25454
rect 36316 25282 36372 25284
rect 36316 25230 36318 25282
rect 36318 25230 36370 25282
rect 36370 25230 36372 25282
rect 36316 25228 36372 25230
rect 36988 24892 37044 24948
rect 36428 24780 36484 24836
rect 37548 25452 37604 25508
rect 37212 24780 37268 24836
rect 37436 25116 37492 25172
rect 35868 23884 35924 23940
rect 36979 24330 37035 24332
rect 36979 24278 36981 24330
rect 36981 24278 37033 24330
rect 37033 24278 37035 24330
rect 36979 24276 37035 24278
rect 37083 24330 37139 24332
rect 37083 24278 37085 24330
rect 37085 24278 37137 24330
rect 37137 24278 37139 24330
rect 37083 24276 37139 24278
rect 37187 24330 37243 24332
rect 37187 24278 37189 24330
rect 37189 24278 37241 24330
rect 37241 24278 37243 24330
rect 37187 24276 37243 24278
rect 38780 25506 38836 25508
rect 38780 25454 38782 25506
rect 38782 25454 38834 25506
rect 38834 25454 38836 25506
rect 38780 25452 38836 25454
rect 37996 25116 38052 25172
rect 36428 23660 36484 23716
rect 38108 23548 38164 23604
rect 34860 21196 34916 21252
rect 34524 20748 34580 20804
rect 33516 20636 33572 20692
rect 34188 20690 34244 20692
rect 34188 20638 34190 20690
rect 34190 20638 34242 20690
rect 34242 20638 34244 20690
rect 34188 20636 34244 20638
rect 35084 20690 35140 20692
rect 35084 20638 35086 20690
rect 35086 20638 35138 20690
rect 35138 20638 35140 20690
rect 35084 20636 35140 20638
rect 34188 20300 34244 20356
rect 33068 20018 33124 20020
rect 33068 19966 33070 20018
rect 33070 19966 33122 20018
rect 33122 19966 33124 20018
rect 33068 19964 33124 19966
rect 34412 19404 34468 19460
rect 33516 19234 33572 19236
rect 33516 19182 33518 19234
rect 33518 19182 33570 19234
rect 33570 19182 33572 19234
rect 33516 19180 33572 19182
rect 33068 17164 33124 17220
rect 33404 18450 33460 18452
rect 33404 18398 33406 18450
rect 33406 18398 33458 18450
rect 33458 18398 33460 18450
rect 33404 18396 33460 18398
rect 33852 19122 33908 19124
rect 33852 19070 33854 19122
rect 33854 19070 33906 19122
rect 33906 19070 33908 19122
rect 33852 19068 33908 19070
rect 33516 17052 33572 17108
rect 33068 16994 33124 16996
rect 33068 16942 33070 16994
rect 33070 16942 33122 16994
rect 33122 16942 33124 16994
rect 33068 16940 33124 16942
rect 33292 16882 33348 16884
rect 33292 16830 33294 16882
rect 33294 16830 33346 16882
rect 33346 16830 33348 16882
rect 33292 16828 33348 16830
rect 33740 17164 33796 17220
rect 33516 16658 33572 16660
rect 33516 16606 33518 16658
rect 33518 16606 33570 16658
rect 33570 16606 33572 16658
rect 33516 16604 33572 16606
rect 34524 18060 34580 18116
rect 34524 17500 34580 17556
rect 34972 19404 35028 19460
rect 35308 21756 35364 21812
rect 35756 23100 35812 23156
rect 35420 21644 35476 21700
rect 35308 19740 35364 19796
rect 34300 17052 34356 17108
rect 34748 18508 34804 18564
rect 33852 16604 33908 16660
rect 33740 16156 33796 16212
rect 34188 15484 34244 15540
rect 33964 15314 34020 15316
rect 33964 15262 33966 15314
rect 33966 15262 34018 15314
rect 34018 15262 34020 15314
rect 33964 15260 34020 15262
rect 34636 16882 34692 16884
rect 34636 16830 34638 16882
rect 34638 16830 34690 16882
rect 34690 16830 34692 16882
rect 34636 16828 34692 16830
rect 35196 18396 35252 18452
rect 35084 18284 35140 18340
rect 34860 18060 34916 18116
rect 34972 17052 35028 17108
rect 34860 16156 34916 16212
rect 35084 15986 35140 15988
rect 35084 15934 35086 15986
rect 35086 15934 35138 15986
rect 35138 15934 35140 15986
rect 35084 15932 35140 15934
rect 32508 14924 32564 14980
rect 33516 14924 33572 14980
rect 32396 14476 32452 14532
rect 33068 13132 33124 13188
rect 32956 12796 33012 12852
rect 32060 12572 32116 12628
rect 32060 11564 32116 11620
rect 32956 12236 33012 12292
rect 34972 15314 35028 15316
rect 34972 15262 34974 15314
rect 34974 15262 35026 15314
rect 35026 15262 35028 15314
rect 34972 15260 35028 15262
rect 35196 15484 35252 15540
rect 34412 14364 34468 14420
rect 34748 13634 34804 13636
rect 34748 13582 34750 13634
rect 34750 13582 34802 13634
rect 34802 13582 34804 13634
rect 34748 13580 34804 13582
rect 34972 13468 35028 13524
rect 33852 12850 33908 12852
rect 33852 12798 33854 12850
rect 33854 12798 33906 12850
rect 33906 12798 33908 12850
rect 33852 12796 33908 12798
rect 35084 12796 35140 12852
rect 34972 12738 35028 12740
rect 34972 12686 34974 12738
rect 34974 12686 35026 12738
rect 35026 12686 35028 12738
rect 34972 12684 35028 12686
rect 34972 12348 35028 12404
rect 33516 12124 33572 12180
rect 34188 12178 34244 12180
rect 34188 12126 34190 12178
rect 34190 12126 34242 12178
rect 34242 12126 34244 12178
rect 34188 12124 34244 12126
rect 33180 11004 33236 11060
rect 35084 12290 35140 12292
rect 35084 12238 35086 12290
rect 35086 12238 35138 12290
rect 35138 12238 35140 12290
rect 35084 12236 35140 12238
rect 35308 12124 35364 12180
rect 36876 23154 36932 23156
rect 36876 23102 36878 23154
rect 36878 23102 36930 23154
rect 36930 23102 36932 23154
rect 36876 23100 36932 23102
rect 36316 23042 36372 23044
rect 36316 22990 36318 23042
rect 36318 22990 36370 23042
rect 36370 22990 36372 23042
rect 36316 22988 36372 22990
rect 35980 22930 36036 22932
rect 35980 22878 35982 22930
rect 35982 22878 36034 22930
rect 36034 22878 36036 22930
rect 35980 22876 36036 22878
rect 37212 22930 37268 22932
rect 37212 22878 37214 22930
rect 37214 22878 37266 22930
rect 37266 22878 37268 22930
rect 37212 22876 37268 22878
rect 36979 22762 37035 22764
rect 36979 22710 36981 22762
rect 36981 22710 37033 22762
rect 37033 22710 37035 22762
rect 36979 22708 37035 22710
rect 37083 22762 37139 22764
rect 37083 22710 37085 22762
rect 37085 22710 37137 22762
rect 37137 22710 37139 22762
rect 37083 22708 37139 22710
rect 37187 22762 37243 22764
rect 37187 22710 37189 22762
rect 37189 22710 37241 22762
rect 37241 22710 37243 22762
rect 37187 22708 37243 22710
rect 36204 22540 36260 22596
rect 36092 20636 36148 20692
rect 36988 22204 37044 22260
rect 36428 21644 36484 21700
rect 37660 23042 37716 23044
rect 37660 22990 37662 23042
rect 37662 22990 37714 23042
rect 37714 22990 37716 23042
rect 37660 22988 37716 22990
rect 38108 22988 38164 23044
rect 37324 21532 37380 21588
rect 37548 22316 37604 22372
rect 40124 26402 40180 26404
rect 40124 26350 40126 26402
rect 40126 26350 40178 26402
rect 40178 26350 40180 26402
rect 40124 26348 40180 26350
rect 39900 26178 39956 26180
rect 39900 26126 39902 26178
rect 39902 26126 39954 26178
rect 39954 26126 39956 26178
rect 39900 26124 39956 26126
rect 40236 26124 40292 26180
rect 46844 26178 46900 26180
rect 46844 26126 46846 26178
rect 46846 26126 46898 26178
rect 46898 26126 46900 26178
rect 46844 26124 46900 26126
rect 41356 25340 41412 25396
rect 40236 25004 40292 25060
rect 39564 24722 39620 24724
rect 39564 24670 39566 24722
rect 39566 24670 39618 24722
rect 39618 24670 39620 24722
rect 39564 24668 39620 24670
rect 39228 23938 39284 23940
rect 39228 23886 39230 23938
rect 39230 23886 39282 23938
rect 39282 23886 39284 23938
rect 39228 23884 39284 23886
rect 39116 23548 39172 23604
rect 38556 22764 38612 22820
rect 38220 22370 38276 22372
rect 38220 22318 38222 22370
rect 38222 22318 38274 22370
rect 38274 22318 38276 22370
rect 38220 22316 38276 22318
rect 39004 22316 39060 22372
rect 38556 22092 38612 22148
rect 36428 20972 36484 21028
rect 36316 20188 36372 20244
rect 36204 19964 36260 20020
rect 35756 19852 35812 19908
rect 35644 19794 35700 19796
rect 35644 19742 35646 19794
rect 35646 19742 35698 19794
rect 35698 19742 35700 19794
rect 35644 19740 35700 19742
rect 36092 19404 36148 19460
rect 35868 19234 35924 19236
rect 35868 19182 35870 19234
rect 35870 19182 35922 19234
rect 35922 19182 35924 19234
rect 35868 19180 35924 19182
rect 35868 18732 35924 18788
rect 35756 18396 35812 18452
rect 36092 18450 36148 18452
rect 36092 18398 36094 18450
rect 36094 18398 36146 18450
rect 36146 18398 36148 18450
rect 36092 18396 36148 18398
rect 35868 18284 35924 18340
rect 35532 17388 35588 17444
rect 35756 17500 35812 17556
rect 36316 17164 36372 17220
rect 36652 19068 36708 19124
rect 36540 18338 36596 18340
rect 36540 18286 36542 18338
rect 36542 18286 36594 18338
rect 36594 18286 36596 18338
rect 36540 18284 36596 18286
rect 36979 21194 37035 21196
rect 36979 21142 36981 21194
rect 36981 21142 37033 21194
rect 37033 21142 37035 21194
rect 36979 21140 37035 21142
rect 37083 21194 37139 21196
rect 37083 21142 37085 21194
rect 37085 21142 37137 21194
rect 37137 21142 37139 21194
rect 37083 21140 37139 21142
rect 37187 21194 37243 21196
rect 37187 21142 37189 21194
rect 37189 21142 37241 21194
rect 37241 21142 37243 21194
rect 37187 21140 37243 21142
rect 36988 20972 37044 21028
rect 37212 20188 37268 20244
rect 36979 19626 37035 19628
rect 36979 19574 36981 19626
rect 36981 19574 37033 19626
rect 37033 19574 37035 19626
rect 36979 19572 37035 19574
rect 37083 19626 37139 19628
rect 37083 19574 37085 19626
rect 37085 19574 37137 19626
rect 37137 19574 37139 19626
rect 37083 19572 37139 19574
rect 37187 19626 37243 19628
rect 37187 19574 37189 19626
rect 37189 19574 37241 19626
rect 37241 19574 37243 19626
rect 37187 19572 37243 19574
rect 37100 18732 37156 18788
rect 37212 19122 37268 19124
rect 37212 19070 37214 19122
rect 37214 19070 37266 19122
rect 37266 19070 37268 19122
rect 37212 19068 37268 19070
rect 37100 18396 37156 18452
rect 36979 18058 37035 18060
rect 36979 18006 36981 18058
rect 36981 18006 37033 18058
rect 37033 18006 37035 18058
rect 36979 18004 37035 18006
rect 37083 18058 37139 18060
rect 37083 18006 37085 18058
rect 37085 18006 37137 18058
rect 37137 18006 37139 18058
rect 37083 18004 37139 18006
rect 37187 18058 37243 18060
rect 37187 18006 37189 18058
rect 37189 18006 37241 18058
rect 37241 18006 37243 18058
rect 37187 18004 37243 18006
rect 37100 17554 37156 17556
rect 37100 17502 37102 17554
rect 37102 17502 37154 17554
rect 37154 17502 37156 17554
rect 37100 17500 37156 17502
rect 36764 16604 36820 16660
rect 36979 16490 37035 16492
rect 36979 16438 36981 16490
rect 36981 16438 37033 16490
rect 37033 16438 37035 16490
rect 36979 16436 37035 16438
rect 37083 16490 37139 16492
rect 37083 16438 37085 16490
rect 37085 16438 37137 16490
rect 37137 16438 37139 16490
rect 37083 16436 37139 16438
rect 37187 16490 37243 16492
rect 37187 16438 37189 16490
rect 37189 16438 37241 16490
rect 37241 16438 37243 16490
rect 37187 16436 37243 16438
rect 36428 16210 36484 16212
rect 36428 16158 36430 16210
rect 36430 16158 36482 16210
rect 36482 16158 36484 16210
rect 36428 16156 36484 16158
rect 36988 16098 37044 16100
rect 36988 16046 36990 16098
rect 36990 16046 37042 16098
rect 37042 16046 37044 16098
rect 36988 16044 37044 16046
rect 36092 15932 36148 15988
rect 36988 15148 37044 15204
rect 35868 15036 35924 15092
rect 35756 14924 35812 14980
rect 37100 15036 37156 15092
rect 38332 21586 38388 21588
rect 38332 21534 38334 21586
rect 38334 21534 38386 21586
rect 38386 21534 38388 21586
rect 38332 21532 38388 21534
rect 38780 20802 38836 20804
rect 38780 20750 38782 20802
rect 38782 20750 38834 20802
rect 38834 20750 38836 20802
rect 38780 20748 38836 20750
rect 38892 20076 38948 20132
rect 37884 20018 37940 20020
rect 37884 19966 37886 20018
rect 37886 19966 37938 20018
rect 37938 19966 37940 20018
rect 37884 19964 37940 19966
rect 38892 19906 38948 19908
rect 38892 19854 38894 19906
rect 38894 19854 38946 19906
rect 38946 19854 38948 19906
rect 38892 19852 38948 19854
rect 37772 19740 37828 19796
rect 37548 17666 37604 17668
rect 37548 17614 37550 17666
rect 37550 17614 37602 17666
rect 37602 17614 37604 17666
rect 37548 17612 37604 17614
rect 38780 18450 38836 18452
rect 38780 18398 38782 18450
rect 38782 18398 38834 18450
rect 38834 18398 38836 18450
rect 38780 18396 38836 18398
rect 39004 17724 39060 17780
rect 39340 23772 39396 23828
rect 41692 24668 41748 24724
rect 41020 23772 41076 23828
rect 39676 23324 39732 23380
rect 40572 23548 40628 23604
rect 40348 23154 40404 23156
rect 40348 23102 40350 23154
rect 40350 23102 40402 23154
rect 40402 23102 40404 23154
rect 40348 23100 40404 23102
rect 39900 23042 39956 23044
rect 39900 22990 39902 23042
rect 39902 22990 39954 23042
rect 39954 22990 39956 23042
rect 39900 22988 39956 22990
rect 39676 22428 39732 22484
rect 40012 22370 40068 22372
rect 40012 22318 40014 22370
rect 40014 22318 40066 22370
rect 40066 22318 40068 22370
rect 40012 22316 40068 22318
rect 40236 21308 40292 21364
rect 39340 19964 39396 20020
rect 39340 19068 39396 19124
rect 40236 20018 40292 20020
rect 40236 19966 40238 20018
rect 40238 19966 40290 20018
rect 40290 19966 40292 20018
rect 40236 19964 40292 19966
rect 40348 19852 40404 19908
rect 40236 19068 40292 19124
rect 39564 17836 39620 17892
rect 39676 18620 39732 18676
rect 37548 17388 37604 17444
rect 37772 16658 37828 16660
rect 37772 16606 37774 16658
rect 37774 16606 37826 16658
rect 37826 16606 37828 16658
rect 37772 16604 37828 16606
rect 37884 16044 37940 16100
rect 37324 15260 37380 15316
rect 36979 14922 37035 14924
rect 36979 14870 36981 14922
rect 36981 14870 37033 14922
rect 37033 14870 37035 14922
rect 36979 14868 37035 14870
rect 37083 14922 37139 14924
rect 37083 14870 37085 14922
rect 37085 14870 37137 14922
rect 37137 14870 37139 14922
rect 37083 14868 37139 14870
rect 37187 14922 37243 14924
rect 37187 14870 37189 14922
rect 37189 14870 37241 14922
rect 37241 14870 37243 14922
rect 37187 14868 37243 14870
rect 35868 14418 35924 14420
rect 35868 14366 35870 14418
rect 35870 14366 35922 14418
rect 35922 14366 35924 14418
rect 35868 14364 35924 14366
rect 36988 14476 37044 14532
rect 35868 13634 35924 13636
rect 35868 13582 35870 13634
rect 35870 13582 35922 13634
rect 35922 13582 35924 13634
rect 35868 13580 35924 13582
rect 35756 13468 35812 13524
rect 35756 12850 35812 12852
rect 35756 12798 35758 12850
rect 35758 12798 35810 12850
rect 35810 12798 35812 12850
rect 35756 12796 35812 12798
rect 35420 12012 35476 12068
rect 35868 12684 35924 12740
rect 36204 14252 36260 14308
rect 36092 13858 36148 13860
rect 36092 13806 36094 13858
rect 36094 13806 36146 13858
rect 36146 13806 36148 13858
rect 36092 13804 36148 13806
rect 35980 12348 36036 12404
rect 33740 9884 33796 9940
rect 32844 9714 32900 9716
rect 32844 9662 32846 9714
rect 32846 9662 32898 9714
rect 32898 9662 32900 9714
rect 32844 9660 32900 9662
rect 29825 9434 29881 9436
rect 29825 9382 29827 9434
rect 29827 9382 29879 9434
rect 29879 9382 29881 9434
rect 29825 9380 29881 9382
rect 29929 9434 29985 9436
rect 29929 9382 29931 9434
rect 29931 9382 29983 9434
rect 29983 9382 29985 9434
rect 29929 9380 29985 9382
rect 30033 9434 30089 9436
rect 30033 9382 30035 9434
rect 30035 9382 30087 9434
rect 30087 9382 30089 9434
rect 30033 9380 30089 9382
rect 29372 8146 29428 8148
rect 29372 8094 29374 8146
rect 29374 8094 29426 8146
rect 29426 8094 29428 8146
rect 29372 8092 29428 8094
rect 27692 7644 27748 7700
rect 28252 7474 28308 7476
rect 28252 7422 28254 7474
rect 28254 7422 28306 7474
rect 28306 7422 28308 7474
rect 28252 7420 28308 7422
rect 27916 7308 27972 7364
rect 28924 7474 28980 7476
rect 28924 7422 28926 7474
rect 28926 7422 28978 7474
rect 28978 7422 28980 7474
rect 28924 7420 28980 7422
rect 27020 5906 27076 5908
rect 27020 5854 27022 5906
rect 27022 5854 27074 5906
rect 27074 5854 27076 5906
rect 27020 5852 27076 5854
rect 27020 5682 27076 5684
rect 27020 5630 27022 5682
rect 27022 5630 27074 5682
rect 27074 5630 27076 5682
rect 27020 5628 27076 5630
rect 27244 5234 27300 5236
rect 27244 5182 27246 5234
rect 27246 5182 27298 5234
rect 27298 5182 27300 5234
rect 27244 5180 27300 5182
rect 27132 4898 27188 4900
rect 27132 4846 27134 4898
rect 27134 4846 27186 4898
rect 27186 4846 27188 4898
rect 27132 4844 27188 4846
rect 26684 4450 26740 4452
rect 26684 4398 26686 4450
rect 26686 4398 26738 4450
rect 26738 4398 26740 4450
rect 26684 4396 26740 4398
rect 27468 4844 27524 4900
rect 26460 4114 26516 4116
rect 26460 4062 26462 4114
rect 26462 4062 26514 4114
rect 26514 4062 26516 4114
rect 26460 4060 26516 4062
rect 27804 5906 27860 5908
rect 27804 5854 27806 5906
rect 27806 5854 27858 5906
rect 27858 5854 27860 5906
rect 27804 5852 27860 5854
rect 28252 6130 28308 6132
rect 28252 6078 28254 6130
rect 28254 6078 28306 6130
rect 28306 6078 28308 6130
rect 28252 6076 28308 6078
rect 28812 6130 28868 6132
rect 28812 6078 28814 6130
rect 28814 6078 28866 6130
rect 28866 6078 28868 6130
rect 28812 6076 28868 6078
rect 29708 8258 29764 8260
rect 29708 8206 29710 8258
rect 29710 8206 29762 8258
rect 29762 8206 29764 8258
rect 29708 8204 29764 8206
rect 29825 7866 29881 7868
rect 29825 7814 29827 7866
rect 29827 7814 29879 7866
rect 29879 7814 29881 7866
rect 29825 7812 29881 7814
rect 29929 7866 29985 7868
rect 29929 7814 29931 7866
rect 29931 7814 29983 7866
rect 29983 7814 29985 7866
rect 29929 7812 29985 7814
rect 30033 7866 30089 7868
rect 30033 7814 30035 7866
rect 30035 7814 30087 7866
rect 30087 7814 30089 7866
rect 30033 7812 30089 7814
rect 29932 7474 29988 7476
rect 29932 7422 29934 7474
rect 29934 7422 29986 7474
rect 29986 7422 29988 7474
rect 29932 7420 29988 7422
rect 30268 7474 30324 7476
rect 30268 7422 30270 7474
rect 30270 7422 30322 7474
rect 30322 7422 30324 7474
rect 30268 7420 30324 7422
rect 29036 5404 29092 5460
rect 29596 6524 29652 6580
rect 29596 6076 29652 6132
rect 28476 5346 28532 5348
rect 28476 5294 28478 5346
rect 28478 5294 28530 5346
rect 28530 5294 28532 5346
rect 28476 5292 28532 5294
rect 31276 8428 31332 8484
rect 31052 8316 31108 8372
rect 31836 8370 31892 8372
rect 31836 8318 31838 8370
rect 31838 8318 31890 8370
rect 31890 8318 31892 8370
rect 31836 8316 31892 8318
rect 33404 8316 33460 8372
rect 31164 8204 31220 8260
rect 32732 8258 32788 8260
rect 32732 8206 32734 8258
rect 32734 8206 32786 8258
rect 32786 8206 32788 8258
rect 32732 8204 32788 8206
rect 36428 12684 36484 12740
rect 35196 11116 35252 11172
rect 36316 11116 36372 11172
rect 35196 8764 35252 8820
rect 30604 6748 30660 6804
rect 30828 6860 30884 6916
rect 29820 6636 29876 6692
rect 29825 6298 29881 6300
rect 29825 6246 29827 6298
rect 29827 6246 29879 6298
rect 29879 6246 29881 6298
rect 29825 6244 29881 6246
rect 29929 6298 29985 6300
rect 29929 6246 29931 6298
rect 29931 6246 29983 6298
rect 29983 6246 29985 6298
rect 29929 6244 29985 6246
rect 30033 6298 30089 6300
rect 30033 6246 30035 6298
rect 30035 6246 30087 6298
rect 30087 6246 30089 6298
rect 30033 6244 30089 6246
rect 29708 5292 29764 5348
rect 30604 5404 30660 5460
rect 32508 8146 32564 8148
rect 32508 8094 32510 8146
rect 32510 8094 32562 8146
rect 32562 8094 32564 8146
rect 32508 8092 32564 8094
rect 33292 8092 33348 8148
rect 33068 8034 33124 8036
rect 33068 7982 33070 8034
rect 33070 7982 33122 8034
rect 33122 7982 33124 8034
rect 33068 7980 33124 7982
rect 32172 7420 32228 7476
rect 31612 6972 31668 7028
rect 33068 7196 33124 7252
rect 31948 6636 32004 6692
rect 32396 6466 32452 6468
rect 32396 6414 32398 6466
rect 32398 6414 32450 6466
rect 32450 6414 32452 6466
rect 32396 6412 32452 6414
rect 31500 5628 31556 5684
rect 28700 4508 28756 4564
rect 28588 4338 28644 4340
rect 28588 4286 28590 4338
rect 28590 4286 28642 4338
rect 28642 4286 28644 4338
rect 28588 4284 28644 4286
rect 28364 4172 28420 4228
rect 30940 5404 30996 5460
rect 29825 4730 29881 4732
rect 29825 4678 29827 4730
rect 29827 4678 29879 4730
rect 29879 4678 29881 4730
rect 29825 4676 29881 4678
rect 29929 4730 29985 4732
rect 29929 4678 29931 4730
rect 29931 4678 29983 4730
rect 29983 4678 29985 4730
rect 29929 4676 29985 4678
rect 30033 4730 30089 4732
rect 30033 4678 30035 4730
rect 30035 4678 30087 4730
rect 30087 4678 30089 4730
rect 30033 4676 30089 4678
rect 29372 4396 29428 4452
rect 32172 5682 32228 5684
rect 32172 5630 32174 5682
rect 32174 5630 32226 5682
rect 32226 5630 32228 5682
rect 32172 5628 32228 5630
rect 32172 5068 32228 5124
rect 32844 6466 32900 6468
rect 32844 6414 32846 6466
rect 32846 6414 32898 6466
rect 32898 6414 32900 6466
rect 32844 6412 32900 6414
rect 33628 8146 33684 8148
rect 33628 8094 33630 8146
rect 33630 8094 33682 8146
rect 33682 8094 33684 8146
rect 33628 8092 33684 8094
rect 36979 13354 37035 13356
rect 36979 13302 36981 13354
rect 36981 13302 37033 13354
rect 37033 13302 37035 13354
rect 36979 13300 37035 13302
rect 37083 13354 37139 13356
rect 37083 13302 37085 13354
rect 37085 13302 37137 13354
rect 37137 13302 37139 13354
rect 37083 13300 37139 13302
rect 37187 13354 37243 13356
rect 37187 13302 37189 13354
rect 37189 13302 37241 13354
rect 37241 13302 37243 13354
rect 37187 13300 37243 13302
rect 37884 14476 37940 14532
rect 37548 14140 37604 14196
rect 38332 14364 38388 14420
rect 38220 14140 38276 14196
rect 37884 13804 37940 13860
rect 37996 13580 38052 13636
rect 37436 13468 37492 13524
rect 37772 12962 37828 12964
rect 37772 12910 37774 12962
rect 37774 12910 37826 12962
rect 37826 12910 37828 12962
rect 37772 12908 37828 12910
rect 37660 12460 37716 12516
rect 41244 23154 41300 23156
rect 41244 23102 41246 23154
rect 41246 23102 41298 23154
rect 41298 23102 41300 23154
rect 41244 23100 41300 23102
rect 41020 22764 41076 22820
rect 41468 22482 41524 22484
rect 41468 22430 41470 22482
rect 41470 22430 41522 22482
rect 41522 22430 41524 22482
rect 41468 22428 41524 22430
rect 41356 22092 41412 22148
rect 42700 25394 42756 25396
rect 42700 25342 42702 25394
rect 42702 25342 42754 25394
rect 42754 25342 42756 25394
rect 42700 25340 42756 25342
rect 42252 24610 42308 24612
rect 42252 24558 42254 24610
rect 42254 24558 42306 24610
rect 42306 24558 42308 24610
rect 42252 24556 42308 24558
rect 42140 23772 42196 23828
rect 42028 23100 42084 23156
rect 42252 23154 42308 23156
rect 42252 23102 42254 23154
rect 42254 23102 42306 23154
rect 42306 23102 42308 23154
rect 42252 23100 42308 23102
rect 42700 24722 42756 24724
rect 42700 24670 42702 24722
rect 42702 24670 42754 24722
rect 42754 24670 42756 24722
rect 42700 24668 42756 24670
rect 48076 26178 48132 26180
rect 48076 26126 48078 26178
rect 48078 26126 48130 26178
rect 48130 26126 48132 26178
rect 48076 26124 48132 26126
rect 48636 26124 48692 26180
rect 47628 25676 47684 25732
rect 47516 25564 47572 25620
rect 44492 25340 44548 25396
rect 42924 24610 42980 24612
rect 42924 24558 42926 24610
rect 42926 24558 42978 24610
rect 42978 24558 42980 24610
rect 42924 24556 42980 24558
rect 42924 23154 42980 23156
rect 42924 23102 42926 23154
rect 42926 23102 42978 23154
rect 42978 23102 42980 23154
rect 42924 23100 42980 23102
rect 44132 25114 44188 25116
rect 44132 25062 44134 25114
rect 44134 25062 44186 25114
rect 44186 25062 44188 25114
rect 44132 25060 44188 25062
rect 44236 25114 44292 25116
rect 44236 25062 44238 25114
rect 44238 25062 44290 25114
rect 44290 25062 44292 25114
rect 44236 25060 44292 25062
rect 44340 25114 44396 25116
rect 44340 25062 44342 25114
rect 44342 25062 44394 25114
rect 44394 25062 44396 25114
rect 44340 25060 44396 25062
rect 43260 24556 43316 24612
rect 44716 25228 44772 25284
rect 45276 25340 45332 25396
rect 45164 25228 45220 25284
rect 45948 24722 46004 24724
rect 45948 24670 45950 24722
rect 45950 24670 46002 24722
rect 46002 24670 46004 24722
rect 45948 24668 46004 24670
rect 46508 24668 46564 24724
rect 47852 25340 47908 25396
rect 48188 25282 48244 25284
rect 48188 25230 48190 25282
rect 48190 25230 48242 25282
rect 48242 25230 48244 25282
rect 48188 25228 48244 25230
rect 48972 25228 49028 25284
rect 46844 23938 46900 23940
rect 46844 23886 46846 23938
rect 46846 23886 46898 23938
rect 46898 23886 46900 23938
rect 46844 23884 46900 23886
rect 44492 23772 44548 23828
rect 43260 23548 43316 23604
rect 44132 23546 44188 23548
rect 44132 23494 44134 23546
rect 44134 23494 44186 23546
rect 44186 23494 44188 23546
rect 44132 23492 44188 23494
rect 44236 23546 44292 23548
rect 44236 23494 44238 23546
rect 44238 23494 44290 23546
rect 44290 23494 44292 23546
rect 44236 23492 44292 23494
rect 44340 23546 44396 23548
rect 44340 23494 44342 23546
rect 44342 23494 44394 23546
rect 44394 23494 44396 23546
rect 44340 23492 44396 23494
rect 43596 22988 43652 23044
rect 42364 22092 42420 22148
rect 42924 22092 42980 22148
rect 40460 18620 40516 18676
rect 40348 18338 40404 18340
rect 40348 18286 40350 18338
rect 40350 18286 40402 18338
rect 40402 18286 40404 18338
rect 40348 18284 40404 18286
rect 40348 17724 40404 17780
rect 39228 16770 39284 16772
rect 39228 16718 39230 16770
rect 39230 16718 39282 16770
rect 39282 16718 39284 16770
rect 39228 16716 39284 16718
rect 38780 16098 38836 16100
rect 38780 16046 38782 16098
rect 38782 16046 38834 16098
rect 38834 16046 38836 16098
rect 38780 16044 38836 16046
rect 39340 15202 39396 15204
rect 39340 15150 39342 15202
rect 39342 15150 39394 15202
rect 39394 15150 39396 15202
rect 39340 15148 39396 15150
rect 40460 17106 40516 17108
rect 40460 17054 40462 17106
rect 40462 17054 40514 17106
rect 40514 17054 40516 17106
rect 40460 17052 40516 17054
rect 40236 15484 40292 15540
rect 40012 15148 40068 15204
rect 42028 21308 42084 21364
rect 41804 20636 41860 20692
rect 41132 19068 41188 19124
rect 41468 18674 41524 18676
rect 41468 18622 41470 18674
rect 41470 18622 41522 18674
rect 41522 18622 41524 18674
rect 41468 18620 41524 18622
rect 41244 18562 41300 18564
rect 41244 18510 41246 18562
rect 41246 18510 41298 18562
rect 41298 18510 41300 18562
rect 41244 18508 41300 18510
rect 41020 17724 41076 17780
rect 41244 18060 41300 18116
rect 41692 19180 41748 19236
rect 42140 21026 42196 21028
rect 42140 20974 42142 21026
rect 42142 20974 42194 21026
rect 42194 20974 42196 21026
rect 42140 20972 42196 20974
rect 42028 20748 42084 20804
rect 42364 20524 42420 20580
rect 42364 20188 42420 20244
rect 42028 20018 42084 20020
rect 42028 19966 42030 20018
rect 42030 19966 42082 20018
rect 42082 19966 42084 20018
rect 42028 19964 42084 19966
rect 42812 19964 42868 20020
rect 42364 19740 42420 19796
rect 42924 19852 42980 19908
rect 41916 19068 41972 19124
rect 43596 21532 43652 21588
rect 43260 19906 43316 19908
rect 43260 19854 43262 19906
rect 43262 19854 43314 19906
rect 43314 19854 43316 19906
rect 43260 19852 43316 19854
rect 44268 22482 44324 22484
rect 44268 22430 44270 22482
rect 44270 22430 44322 22482
rect 44322 22430 44324 22482
rect 44268 22428 44324 22430
rect 43708 20972 43764 21028
rect 43820 20188 43876 20244
rect 44828 22316 44884 22372
rect 44044 22092 44100 22148
rect 44132 21978 44188 21980
rect 44132 21926 44134 21978
rect 44134 21926 44186 21978
rect 44186 21926 44188 21978
rect 44132 21924 44188 21926
rect 44236 21978 44292 21980
rect 44236 21926 44238 21978
rect 44238 21926 44290 21978
rect 44290 21926 44292 21978
rect 44236 21924 44292 21926
rect 44340 21978 44396 21980
rect 44340 21926 44342 21978
rect 44342 21926 44394 21978
rect 44394 21926 44396 21978
rect 44340 21924 44396 21926
rect 44044 21420 44100 21476
rect 44492 20748 44548 20804
rect 44044 20690 44100 20692
rect 44044 20638 44046 20690
rect 44046 20638 44098 20690
rect 44098 20638 44100 20690
rect 44044 20636 44100 20638
rect 44132 20410 44188 20412
rect 44132 20358 44134 20410
rect 44134 20358 44186 20410
rect 44186 20358 44188 20410
rect 44132 20356 44188 20358
rect 44236 20410 44292 20412
rect 44236 20358 44238 20410
rect 44238 20358 44290 20410
rect 44290 20358 44292 20410
rect 44236 20356 44292 20358
rect 44340 20410 44396 20412
rect 44340 20358 44342 20410
rect 44342 20358 44394 20410
rect 44394 20358 44396 20410
rect 44340 20356 44396 20358
rect 44380 20188 44436 20244
rect 43932 19458 43988 19460
rect 43932 19406 43934 19458
rect 43934 19406 43986 19458
rect 43986 19406 43988 19458
rect 43932 19404 43988 19406
rect 41804 18284 41860 18340
rect 42140 18172 42196 18228
rect 41580 18060 41636 18116
rect 42252 17890 42308 17892
rect 42252 17838 42254 17890
rect 42254 17838 42306 17890
rect 42306 17838 42308 17890
rect 42252 17836 42308 17838
rect 41692 17724 41748 17780
rect 41244 17052 41300 17108
rect 42252 17388 42308 17444
rect 41580 16828 41636 16884
rect 42140 17106 42196 17108
rect 42140 17054 42142 17106
rect 42142 17054 42194 17106
rect 42194 17054 42196 17106
rect 42140 17052 42196 17054
rect 42812 18508 42868 18564
rect 44156 19180 44212 19236
rect 44132 18842 44188 18844
rect 44132 18790 44134 18842
rect 44134 18790 44186 18842
rect 44186 18790 44188 18842
rect 44132 18788 44188 18790
rect 44236 18842 44292 18844
rect 44236 18790 44238 18842
rect 44238 18790 44290 18842
rect 44290 18790 44292 18842
rect 44236 18788 44292 18790
rect 44340 18842 44396 18844
rect 44340 18790 44342 18842
rect 44342 18790 44394 18842
rect 44394 18790 44396 18842
rect 44340 18788 44396 18790
rect 42924 18450 42980 18452
rect 42924 18398 42926 18450
rect 42926 18398 42978 18450
rect 42978 18398 42980 18450
rect 42924 18396 42980 18398
rect 42812 17836 42868 17892
rect 42476 17276 42532 17332
rect 43260 18060 43316 18116
rect 43148 17442 43204 17444
rect 43148 17390 43150 17442
rect 43150 17390 43202 17442
rect 43202 17390 43204 17442
rect 43148 17388 43204 17390
rect 42588 16828 42644 16884
rect 40908 15260 40964 15316
rect 41244 15260 41300 15316
rect 39564 14642 39620 14644
rect 39564 14590 39566 14642
rect 39566 14590 39618 14642
rect 39618 14590 39620 14642
rect 39564 14588 39620 14590
rect 39228 14418 39284 14420
rect 39228 14366 39230 14418
rect 39230 14366 39282 14418
rect 39282 14366 39284 14418
rect 39228 14364 39284 14366
rect 38444 13580 38500 13636
rect 38668 14140 38724 14196
rect 39228 13468 39284 13524
rect 38668 12460 38724 12516
rect 38332 12012 38388 12068
rect 36979 11786 37035 11788
rect 36764 11676 36820 11732
rect 36979 11734 36981 11786
rect 36981 11734 37033 11786
rect 37033 11734 37035 11786
rect 36979 11732 37035 11734
rect 37083 11786 37139 11788
rect 37083 11734 37085 11786
rect 37085 11734 37137 11786
rect 37137 11734 37139 11786
rect 37083 11732 37139 11734
rect 37187 11786 37243 11788
rect 37187 11734 37189 11786
rect 37189 11734 37241 11786
rect 37241 11734 37243 11786
rect 37187 11732 37243 11734
rect 36764 11452 36820 11508
rect 38220 11170 38276 11172
rect 38220 11118 38222 11170
rect 38222 11118 38274 11170
rect 38274 11118 38276 11170
rect 38220 11116 38276 11118
rect 37772 10780 37828 10836
rect 37660 10386 37716 10388
rect 37660 10334 37662 10386
rect 37662 10334 37714 10386
rect 37714 10334 37716 10386
rect 37660 10332 37716 10334
rect 36979 10218 37035 10220
rect 36979 10166 36981 10218
rect 36981 10166 37033 10218
rect 37033 10166 37035 10218
rect 36979 10164 37035 10166
rect 37083 10218 37139 10220
rect 37083 10166 37085 10218
rect 37085 10166 37137 10218
rect 37137 10166 37139 10218
rect 37083 10164 37139 10166
rect 37187 10218 37243 10220
rect 37187 10166 37189 10218
rect 37189 10166 37241 10218
rect 37241 10166 37243 10218
rect 37187 10164 37243 10166
rect 38332 10834 38388 10836
rect 38332 10782 38334 10834
rect 38334 10782 38386 10834
rect 38386 10782 38388 10834
rect 38332 10780 38388 10782
rect 39900 14364 39956 14420
rect 39452 14140 39508 14196
rect 39564 13804 39620 13860
rect 39564 13468 39620 13524
rect 40124 13580 40180 13636
rect 40348 12962 40404 12964
rect 40348 12910 40350 12962
rect 40350 12910 40402 12962
rect 40402 12910 40404 12962
rect 40348 12908 40404 12910
rect 39900 11004 39956 11060
rect 40572 14588 40628 14644
rect 41020 13522 41076 13524
rect 41020 13470 41022 13522
rect 41022 13470 41074 13522
rect 41074 13470 41076 13522
rect 41020 13468 41076 13470
rect 40236 11116 40292 11172
rect 40684 11170 40740 11172
rect 40684 11118 40686 11170
rect 40686 11118 40738 11170
rect 40738 11118 40740 11170
rect 40684 11116 40740 11118
rect 36428 9884 36484 9940
rect 36428 9548 36484 9604
rect 37100 9548 37156 9604
rect 36979 8650 37035 8652
rect 36979 8598 36981 8650
rect 36981 8598 37033 8650
rect 37033 8598 37035 8650
rect 36979 8596 37035 8598
rect 37083 8650 37139 8652
rect 37083 8598 37085 8650
rect 37085 8598 37137 8650
rect 37137 8598 37139 8650
rect 37083 8596 37139 8598
rect 37187 8650 37243 8652
rect 37187 8598 37189 8650
rect 37189 8598 37241 8650
rect 37241 8598 37243 8650
rect 37187 8596 37243 8598
rect 37548 8428 37604 8484
rect 36092 8316 36148 8372
rect 34076 8092 34132 8148
rect 34972 8146 35028 8148
rect 34972 8094 34974 8146
rect 34974 8094 35026 8146
rect 35026 8094 35028 8146
rect 34972 8092 35028 8094
rect 35532 8146 35588 8148
rect 35532 8094 35534 8146
rect 35534 8094 35586 8146
rect 35586 8094 35588 8146
rect 35532 8092 35588 8094
rect 34524 7980 34580 8036
rect 34188 7586 34244 7588
rect 34188 7534 34190 7586
rect 34190 7534 34242 7586
rect 34242 7534 34244 7586
rect 34188 7532 34244 7534
rect 33964 7250 34020 7252
rect 33964 7198 33966 7250
rect 33966 7198 34018 7250
rect 34018 7198 34020 7250
rect 33964 7196 34020 7198
rect 33740 6636 33796 6692
rect 31164 4284 31220 4340
rect 28924 4172 28980 4228
rect 25676 3666 25732 3668
rect 25676 3614 25678 3666
rect 25678 3614 25730 3666
rect 25730 3614 25732 3666
rect 25676 3612 25732 3614
rect 31948 3948 32004 4004
rect 27356 3612 27412 3668
rect 35084 8034 35140 8036
rect 35084 7982 35086 8034
rect 35086 7982 35138 8034
rect 35138 7982 35140 8034
rect 35084 7980 35140 7982
rect 35420 7980 35476 8036
rect 34748 7474 34804 7476
rect 34748 7422 34750 7474
rect 34750 7422 34802 7474
rect 34802 7422 34804 7474
rect 34748 7420 34804 7422
rect 34636 6690 34692 6692
rect 34636 6638 34638 6690
rect 34638 6638 34690 6690
rect 34690 6638 34692 6690
rect 34636 6636 34692 6638
rect 35644 7532 35700 7588
rect 32284 4338 32340 4340
rect 32284 4286 32286 4338
rect 32286 4286 32338 4338
rect 32338 4286 32340 4338
rect 32284 4284 32340 4286
rect 25452 3500 25508 3556
rect 33404 5180 33460 5236
rect 34412 5234 34468 5236
rect 34412 5182 34414 5234
rect 34414 5182 34466 5234
rect 34466 5182 34468 5234
rect 34412 5180 34468 5182
rect 35196 5906 35252 5908
rect 35196 5854 35198 5906
rect 35198 5854 35250 5906
rect 35250 5854 35252 5906
rect 35196 5852 35252 5854
rect 35084 5794 35140 5796
rect 35084 5742 35086 5794
rect 35086 5742 35138 5794
rect 35138 5742 35140 5794
rect 35084 5740 35140 5742
rect 35420 6636 35476 6692
rect 35756 5852 35812 5908
rect 35868 5628 35924 5684
rect 35420 4732 35476 4788
rect 36979 7082 37035 7084
rect 36979 7030 36981 7082
rect 36981 7030 37033 7082
rect 37033 7030 37035 7082
rect 36979 7028 37035 7030
rect 37083 7082 37139 7084
rect 37083 7030 37085 7082
rect 37085 7030 37137 7082
rect 37137 7030 37139 7082
rect 37083 7028 37139 7030
rect 37187 7082 37243 7084
rect 37187 7030 37189 7082
rect 37189 7030 37241 7082
rect 37241 7030 37243 7082
rect 37187 7028 37243 7030
rect 36092 4732 36148 4788
rect 36316 6636 36372 6692
rect 36988 6130 37044 6132
rect 36988 6078 36990 6130
rect 36990 6078 37042 6130
rect 37042 6078 37044 6130
rect 36988 6076 37044 6078
rect 36979 5514 37035 5516
rect 36979 5462 36981 5514
rect 36981 5462 37033 5514
rect 37033 5462 37035 5514
rect 36979 5460 37035 5462
rect 37083 5514 37139 5516
rect 37083 5462 37085 5514
rect 37085 5462 37137 5514
rect 37137 5462 37139 5514
rect 37083 5460 37139 5462
rect 37187 5514 37243 5516
rect 37187 5462 37189 5514
rect 37189 5462 37241 5514
rect 37241 5462 37243 5514
rect 37187 5460 37243 5462
rect 36876 4956 36932 5012
rect 33068 4338 33124 4340
rect 33068 4286 33070 4338
rect 33070 4286 33122 4338
rect 33122 4286 33124 4338
rect 33068 4284 33124 4286
rect 33292 3948 33348 4004
rect 38444 9938 38500 9940
rect 38444 9886 38446 9938
rect 38446 9886 38498 9938
rect 38498 9886 38500 9938
rect 38444 9884 38500 9886
rect 37772 9772 37828 9828
rect 38108 9660 38164 9716
rect 38108 8204 38164 8260
rect 37548 6130 37604 6132
rect 37548 6078 37550 6130
rect 37550 6078 37602 6130
rect 37602 6078 37604 6130
rect 37548 6076 37604 6078
rect 37884 5906 37940 5908
rect 37884 5854 37886 5906
rect 37886 5854 37938 5906
rect 37938 5854 37940 5906
rect 37884 5852 37940 5854
rect 37660 5404 37716 5460
rect 37436 4620 37492 4676
rect 36979 3946 37035 3948
rect 36979 3894 36981 3946
rect 36981 3894 37033 3946
rect 37033 3894 37035 3946
rect 36979 3892 37035 3894
rect 37083 3946 37139 3948
rect 37083 3894 37085 3946
rect 37085 3894 37137 3946
rect 37137 3894 37139 3946
rect 37083 3892 37139 3894
rect 37187 3946 37243 3948
rect 37187 3894 37189 3946
rect 37189 3894 37241 3946
rect 37241 3894 37243 3946
rect 37187 3892 37243 3894
rect 37548 3554 37604 3556
rect 37548 3502 37550 3554
rect 37550 3502 37602 3554
rect 37602 3502 37604 3554
rect 37548 3500 37604 3502
rect 25788 3442 25844 3444
rect 25788 3390 25790 3442
rect 25790 3390 25842 3442
rect 25842 3390 25844 3442
rect 25788 3388 25844 3390
rect 38332 9714 38388 9716
rect 38332 9662 38334 9714
rect 38334 9662 38386 9714
rect 38386 9662 38388 9714
rect 38332 9660 38388 9662
rect 39340 9714 39396 9716
rect 39340 9662 39342 9714
rect 39342 9662 39394 9714
rect 39394 9662 39396 9714
rect 39340 9660 39396 9662
rect 39452 9266 39508 9268
rect 39452 9214 39454 9266
rect 39454 9214 39506 9266
rect 39506 9214 39508 9266
rect 39452 9212 39508 9214
rect 39228 8204 39284 8260
rect 39004 6578 39060 6580
rect 39004 6526 39006 6578
rect 39006 6526 39058 6578
rect 39058 6526 39060 6578
rect 39004 6524 39060 6526
rect 39788 9884 39844 9940
rect 40124 10780 40180 10836
rect 41244 13916 41300 13972
rect 42140 15538 42196 15540
rect 42140 15486 42142 15538
rect 42142 15486 42194 15538
rect 42194 15486 42196 15538
rect 42140 15484 42196 15486
rect 44132 17274 44188 17276
rect 44132 17222 44134 17274
rect 44134 17222 44186 17274
rect 44186 17222 44188 17274
rect 44132 17220 44188 17222
rect 44236 17274 44292 17276
rect 44236 17222 44238 17274
rect 44238 17222 44290 17274
rect 44290 17222 44292 17274
rect 44236 17220 44292 17222
rect 44340 17274 44396 17276
rect 44340 17222 44342 17274
rect 44342 17222 44394 17274
rect 44394 17222 44396 17274
rect 44340 17220 44396 17222
rect 43708 16716 43764 16772
rect 45276 22204 45332 22260
rect 45948 21644 46004 21700
rect 44940 20524 44996 20580
rect 46060 20802 46116 20804
rect 46060 20750 46062 20802
rect 46062 20750 46114 20802
rect 46114 20750 46116 20802
rect 46060 20748 46116 20750
rect 45836 20188 45892 20244
rect 45948 20076 46004 20132
rect 45276 19740 45332 19796
rect 47180 23772 47236 23828
rect 47068 23154 47124 23156
rect 47068 23102 47070 23154
rect 47070 23102 47122 23154
rect 47122 23102 47124 23154
rect 47068 23100 47124 23102
rect 46508 22428 46564 22484
rect 46508 21868 46564 21924
rect 46956 22540 47012 22596
rect 46284 20018 46340 20020
rect 46284 19966 46286 20018
rect 46286 19966 46338 20018
rect 46338 19966 46340 20018
rect 46284 19964 46340 19966
rect 46620 21420 46676 21476
rect 46172 19794 46228 19796
rect 46172 19742 46174 19794
rect 46174 19742 46226 19794
rect 46226 19742 46228 19794
rect 46172 19740 46228 19742
rect 45276 19180 45332 19236
rect 44604 18284 44660 18340
rect 44716 17612 44772 17668
rect 45164 19010 45220 19012
rect 45164 18958 45166 19010
rect 45166 18958 45218 19010
rect 45218 18958 45220 19010
rect 45164 18956 45220 18958
rect 43932 16098 43988 16100
rect 43932 16046 43934 16098
rect 43934 16046 43986 16098
rect 43986 16046 43988 16098
rect 43932 16044 43988 16046
rect 43820 15874 43876 15876
rect 43820 15822 43822 15874
rect 43822 15822 43874 15874
rect 43874 15822 43876 15874
rect 43820 15820 43876 15822
rect 46060 19628 46116 19684
rect 46508 19516 46564 19572
rect 45276 18060 45332 18116
rect 46732 20802 46788 20804
rect 46732 20750 46734 20802
rect 46734 20750 46786 20802
rect 46786 20750 46788 20802
rect 46732 20748 46788 20750
rect 47068 22370 47124 22372
rect 47068 22318 47070 22370
rect 47070 22318 47122 22370
rect 47122 22318 47124 22370
rect 47068 22316 47124 22318
rect 47292 22316 47348 22372
rect 48188 24610 48244 24612
rect 48188 24558 48190 24610
rect 48190 24558 48242 24610
rect 48242 24558 48244 24610
rect 48188 24556 48244 24558
rect 47964 22258 48020 22260
rect 47964 22206 47966 22258
rect 47966 22206 48018 22258
rect 48018 22206 48020 22258
rect 47964 22204 48020 22206
rect 47740 22092 47796 22148
rect 47180 20972 47236 21028
rect 47404 21420 47460 21476
rect 46844 19628 46900 19684
rect 47068 20130 47124 20132
rect 47068 20078 47070 20130
rect 47070 20078 47122 20130
rect 47122 20078 47124 20130
rect 47068 20076 47124 20078
rect 46956 19964 47012 20020
rect 46732 19404 46788 19460
rect 46732 18450 46788 18452
rect 46732 18398 46734 18450
rect 46734 18398 46786 18450
rect 46786 18398 46788 18450
rect 46732 18396 46788 18398
rect 46956 19180 47012 19236
rect 47180 19852 47236 19908
rect 46844 18284 46900 18340
rect 46284 17666 46340 17668
rect 46284 17614 46286 17666
rect 46286 17614 46338 17666
rect 46338 17614 46340 17666
rect 46284 17612 46340 17614
rect 45388 17106 45444 17108
rect 45388 17054 45390 17106
rect 45390 17054 45442 17106
rect 45442 17054 45444 17106
rect 45388 17052 45444 17054
rect 45052 16098 45108 16100
rect 45052 16046 45054 16098
rect 45054 16046 45106 16098
rect 45106 16046 45108 16098
rect 45052 16044 45108 16046
rect 45836 15932 45892 15988
rect 44132 15706 44188 15708
rect 44132 15654 44134 15706
rect 44134 15654 44186 15706
rect 44186 15654 44188 15706
rect 44132 15652 44188 15654
rect 44236 15706 44292 15708
rect 44236 15654 44238 15706
rect 44238 15654 44290 15706
rect 44290 15654 44292 15706
rect 44236 15652 44292 15654
rect 44340 15706 44396 15708
rect 44340 15654 44342 15706
rect 44342 15654 44394 15706
rect 44394 15654 44396 15706
rect 44340 15652 44396 15654
rect 44604 15538 44660 15540
rect 44604 15486 44606 15538
rect 44606 15486 44658 15538
rect 44658 15486 44660 15538
rect 44604 15484 44660 15486
rect 45724 15820 45780 15876
rect 41580 15260 41636 15316
rect 42364 15314 42420 15316
rect 42364 15262 42366 15314
rect 42366 15262 42418 15314
rect 42418 15262 42420 15314
rect 42364 15260 42420 15262
rect 41580 13858 41636 13860
rect 41580 13806 41582 13858
rect 41582 13806 41634 13858
rect 41634 13806 41636 13858
rect 41580 13804 41636 13806
rect 41692 13916 41748 13972
rect 41244 13580 41300 13636
rect 40348 10108 40404 10164
rect 40124 9884 40180 9940
rect 40012 9212 40068 9268
rect 41244 9996 41300 10052
rect 40908 9660 40964 9716
rect 40460 9100 40516 9156
rect 40236 8876 40292 8932
rect 40124 7474 40180 7476
rect 40124 7422 40126 7474
rect 40126 7422 40178 7474
rect 40178 7422 40180 7474
rect 40124 7420 40180 7422
rect 40124 6636 40180 6692
rect 38332 5404 38388 5460
rect 38444 5180 38500 5236
rect 38556 6188 38612 6244
rect 39004 6188 39060 6244
rect 38220 4956 38276 5012
rect 38668 5068 38724 5124
rect 39900 6130 39956 6132
rect 39900 6078 39902 6130
rect 39902 6078 39954 6130
rect 39954 6078 39956 6130
rect 39900 6076 39956 6078
rect 39452 5852 39508 5908
rect 39228 5180 39284 5236
rect 39116 4898 39172 4900
rect 39116 4846 39118 4898
rect 39118 4846 39170 4898
rect 39170 4846 39172 4898
rect 39116 4844 39172 4846
rect 40572 8428 40628 8484
rect 40908 8988 40964 9044
rect 40796 8428 40852 8484
rect 42028 13746 42084 13748
rect 42028 13694 42030 13746
rect 42030 13694 42082 13746
rect 42082 13694 42084 13746
rect 42028 13692 42084 13694
rect 42252 13468 42308 13524
rect 41692 11004 41748 11060
rect 41580 9154 41636 9156
rect 41580 9102 41582 9154
rect 41582 9102 41634 9154
rect 41634 9102 41636 9154
rect 41580 9100 41636 9102
rect 41020 8316 41076 8372
rect 41916 10610 41972 10612
rect 41916 10558 41918 10610
rect 41918 10558 41970 10610
rect 41970 10558 41972 10610
rect 41916 10556 41972 10558
rect 41692 8316 41748 8372
rect 42028 9100 42084 9156
rect 42140 9996 42196 10052
rect 41804 8258 41860 8260
rect 41804 8206 41806 8258
rect 41806 8206 41858 8258
rect 41858 8206 41860 8258
rect 41804 8204 41860 8206
rect 42700 14700 42756 14756
rect 45388 15538 45444 15540
rect 45388 15486 45390 15538
rect 45390 15486 45442 15538
rect 45442 15486 45444 15538
rect 45388 15484 45444 15486
rect 47404 20524 47460 20580
rect 47628 21756 47684 21812
rect 47404 19516 47460 19572
rect 47516 20130 47572 20132
rect 47516 20078 47518 20130
rect 47518 20078 47570 20130
rect 47570 20078 47572 20130
rect 47516 20076 47572 20078
rect 48636 23884 48692 23940
rect 50316 26514 50372 26516
rect 50316 26462 50318 26514
rect 50318 26462 50370 26514
rect 50370 26462 50372 26514
rect 50316 26460 50372 26462
rect 52220 26514 52276 26516
rect 52220 26462 52222 26514
rect 52222 26462 52274 26514
rect 52274 26462 52276 26514
rect 52220 26460 52276 26462
rect 58439 26682 58495 26684
rect 58439 26630 58441 26682
rect 58441 26630 58493 26682
rect 58493 26630 58495 26682
rect 58439 26628 58495 26630
rect 58543 26682 58599 26684
rect 58543 26630 58545 26682
rect 58545 26630 58597 26682
rect 58597 26630 58599 26682
rect 58543 26628 58599 26630
rect 58647 26682 58703 26684
rect 58647 26630 58649 26682
rect 58649 26630 58701 26682
rect 58701 26630 58703 26682
rect 58647 26628 58703 26630
rect 49532 26290 49588 26292
rect 49532 26238 49534 26290
rect 49534 26238 49586 26290
rect 49586 26238 49588 26290
rect 49532 26236 49588 26238
rect 49196 26066 49252 26068
rect 49196 26014 49198 26066
rect 49198 26014 49250 26066
rect 49250 26014 49252 26066
rect 49196 26012 49252 26014
rect 49980 26290 50036 26292
rect 49980 26238 49982 26290
rect 49982 26238 50034 26290
rect 50034 26238 50036 26290
rect 49980 26236 50036 26238
rect 50428 26236 50484 26292
rect 50204 26012 50260 26068
rect 49196 25394 49252 25396
rect 49196 25342 49198 25394
rect 49198 25342 49250 25394
rect 49250 25342 49252 25394
rect 49196 25340 49252 25342
rect 48748 23772 48804 23828
rect 48412 23100 48468 23156
rect 49532 23266 49588 23268
rect 49532 23214 49534 23266
rect 49534 23214 49586 23266
rect 49586 23214 49588 23266
rect 49532 23212 49588 23214
rect 48748 22428 48804 22484
rect 48972 21980 49028 22036
rect 48188 21474 48244 21476
rect 48188 21422 48190 21474
rect 48190 21422 48242 21474
rect 48242 21422 48244 21474
rect 48188 21420 48244 21422
rect 47964 20524 48020 20580
rect 47628 18396 47684 18452
rect 48076 20412 48132 20468
rect 48748 21586 48804 21588
rect 48748 21534 48750 21586
rect 48750 21534 48802 21586
rect 48802 21534 48804 21586
rect 48748 21532 48804 21534
rect 49308 21698 49364 21700
rect 49308 21646 49310 21698
rect 49310 21646 49362 21698
rect 49362 21646 49364 21698
rect 49308 21644 49364 21646
rect 48636 21420 48692 21476
rect 49532 22370 49588 22372
rect 49532 22318 49534 22370
rect 49534 22318 49586 22370
rect 49586 22318 49588 22370
rect 49532 22316 49588 22318
rect 49532 21868 49588 21924
rect 49644 21756 49700 21812
rect 48188 18508 48244 18564
rect 48076 18396 48132 18452
rect 48972 19628 49028 19684
rect 49420 20018 49476 20020
rect 49420 19966 49422 20018
rect 49422 19966 49474 20018
rect 49474 19966 49476 20018
rect 49420 19964 49476 19966
rect 49308 19906 49364 19908
rect 49308 19854 49310 19906
rect 49310 19854 49362 19906
rect 49362 19854 49364 19906
rect 49308 19852 49364 19854
rect 48860 18562 48916 18564
rect 48860 18510 48862 18562
rect 48862 18510 48914 18562
rect 48914 18510 48916 18562
rect 48860 18508 48916 18510
rect 49196 18284 49252 18340
rect 48748 18172 48804 18228
rect 49420 18508 49476 18564
rect 49756 23212 49812 23268
rect 49756 22204 49812 22260
rect 49868 19234 49924 19236
rect 49868 19182 49870 19234
rect 49870 19182 49922 19234
rect 49922 19182 49924 19234
rect 49868 19180 49924 19182
rect 49532 18284 49588 18340
rect 49756 18620 49812 18676
rect 49308 17106 49364 17108
rect 49308 17054 49310 17106
rect 49310 17054 49362 17106
rect 49362 17054 49364 17106
rect 49308 17052 49364 17054
rect 46508 15986 46564 15988
rect 46508 15934 46510 15986
rect 46510 15934 46562 15986
rect 46562 15934 46564 15986
rect 46508 15932 46564 15934
rect 47628 15932 47684 15988
rect 48972 16098 49028 16100
rect 48972 16046 48974 16098
rect 48974 16046 49026 16098
rect 49026 16046 49028 16098
rect 48972 16044 49028 16046
rect 47964 15932 48020 15988
rect 47852 15426 47908 15428
rect 47852 15374 47854 15426
rect 47854 15374 47906 15426
rect 47906 15374 47908 15426
rect 47852 15372 47908 15374
rect 44268 14476 44324 14532
rect 44828 14530 44884 14532
rect 44828 14478 44830 14530
rect 44830 14478 44882 14530
rect 44882 14478 44884 14530
rect 44828 14476 44884 14478
rect 44604 14364 44660 14420
rect 45276 14418 45332 14420
rect 45276 14366 45278 14418
rect 45278 14366 45330 14418
rect 45330 14366 45332 14418
rect 45276 14364 45332 14366
rect 45836 14364 45892 14420
rect 47516 15314 47572 15316
rect 47516 15262 47518 15314
rect 47518 15262 47570 15314
rect 47570 15262 47572 15314
rect 47516 15260 47572 15262
rect 44132 14138 44188 14140
rect 44132 14086 44134 14138
rect 44134 14086 44186 14138
rect 44186 14086 44188 14138
rect 44132 14084 44188 14086
rect 44236 14138 44292 14140
rect 44236 14086 44238 14138
rect 44238 14086 44290 14138
rect 44290 14086 44292 14138
rect 44236 14084 44292 14086
rect 44340 14138 44396 14140
rect 44340 14086 44342 14138
rect 44342 14086 44394 14138
rect 44394 14086 44396 14138
rect 44340 14084 44396 14086
rect 44604 13858 44660 13860
rect 44604 13806 44606 13858
rect 44606 13806 44658 13858
rect 44658 13806 44660 13858
rect 44604 13804 44660 13806
rect 45500 13858 45556 13860
rect 45500 13806 45502 13858
rect 45502 13806 45554 13858
rect 45554 13806 45556 13858
rect 45500 13804 45556 13806
rect 42700 12348 42756 12404
rect 45724 13746 45780 13748
rect 45724 13694 45726 13746
rect 45726 13694 45778 13746
rect 45778 13694 45780 13746
rect 45724 13692 45780 13694
rect 46732 13132 46788 13188
rect 45164 13074 45220 13076
rect 45164 13022 45166 13074
rect 45166 13022 45218 13074
rect 45218 13022 45220 13074
rect 45164 13020 45220 13022
rect 47292 13186 47348 13188
rect 47292 13134 47294 13186
rect 47294 13134 47346 13186
rect 47346 13134 47348 13186
rect 47292 13132 47348 13134
rect 44940 12908 44996 12964
rect 45500 12962 45556 12964
rect 45500 12910 45502 12962
rect 45502 12910 45554 12962
rect 45554 12910 45556 12962
rect 45500 12908 45556 12910
rect 45836 12738 45892 12740
rect 45836 12686 45838 12738
rect 45838 12686 45890 12738
rect 45890 12686 45892 12738
rect 45836 12684 45892 12686
rect 42924 11788 42980 11844
rect 44132 12570 44188 12572
rect 44132 12518 44134 12570
rect 44134 12518 44186 12570
rect 44186 12518 44188 12570
rect 44132 12516 44188 12518
rect 44236 12570 44292 12572
rect 44236 12518 44238 12570
rect 44238 12518 44290 12570
rect 44290 12518 44292 12570
rect 44236 12516 44292 12518
rect 44340 12570 44396 12572
rect 44340 12518 44342 12570
rect 44342 12518 44394 12570
rect 44394 12518 44396 12570
rect 44340 12516 44396 12518
rect 47068 12684 47124 12740
rect 44380 12402 44436 12404
rect 44380 12350 44382 12402
rect 44382 12350 44434 12402
rect 44434 12350 44436 12402
rect 44380 12348 44436 12350
rect 45164 12348 45220 12404
rect 47292 12236 47348 12292
rect 48188 15202 48244 15204
rect 48188 15150 48190 15202
rect 48190 15150 48242 15202
rect 48242 15150 48244 15202
rect 48188 15148 48244 15150
rect 47516 14418 47572 14420
rect 47516 14366 47518 14418
rect 47518 14366 47570 14418
rect 47570 14366 47572 14418
rect 47516 14364 47572 14366
rect 49308 15932 49364 15988
rect 49196 15148 49252 15204
rect 48188 14140 48244 14196
rect 47852 13692 47908 13748
rect 47516 12738 47572 12740
rect 47516 12686 47518 12738
rect 47518 12686 47570 12738
rect 47570 12686 47572 12738
rect 47516 12684 47572 12686
rect 47516 12402 47572 12404
rect 47516 12350 47518 12402
rect 47518 12350 47570 12402
rect 47570 12350 47572 12402
rect 47516 12348 47572 12350
rect 47852 12402 47908 12404
rect 47852 12350 47854 12402
rect 47854 12350 47906 12402
rect 47906 12350 47908 12402
rect 47852 12348 47908 12350
rect 48748 14140 48804 14196
rect 48524 13132 48580 13188
rect 48076 12962 48132 12964
rect 48076 12910 48078 12962
rect 48078 12910 48130 12962
rect 48130 12910 48132 12962
rect 48076 12908 48132 12910
rect 48524 12962 48580 12964
rect 48524 12910 48526 12962
rect 48526 12910 48578 12962
rect 48578 12910 48580 12962
rect 48524 12908 48580 12910
rect 48748 13468 48804 13524
rect 49868 15036 49924 15092
rect 50092 20130 50148 20132
rect 50092 20078 50094 20130
rect 50094 20078 50146 20130
rect 50146 20078 50148 20130
rect 50092 20076 50148 20078
rect 50428 26012 50484 26068
rect 51772 26178 51828 26180
rect 51772 26126 51774 26178
rect 51774 26126 51826 26178
rect 51826 26126 51828 26178
rect 51772 26124 51828 26126
rect 51212 26066 51268 26068
rect 51212 26014 51214 26066
rect 51214 26014 51266 26066
rect 51266 26014 51268 26066
rect 51212 26012 51268 26014
rect 51286 25898 51342 25900
rect 51286 25846 51288 25898
rect 51288 25846 51340 25898
rect 51340 25846 51342 25898
rect 51286 25844 51342 25846
rect 51390 25898 51446 25900
rect 51390 25846 51392 25898
rect 51392 25846 51444 25898
rect 51444 25846 51446 25898
rect 51390 25844 51446 25846
rect 51494 25898 51550 25900
rect 51494 25846 51496 25898
rect 51496 25846 51548 25898
rect 51548 25846 51550 25898
rect 51494 25844 51550 25846
rect 50540 24556 50596 24612
rect 51286 24330 51342 24332
rect 51286 24278 51288 24330
rect 51288 24278 51340 24330
rect 51340 24278 51342 24330
rect 51286 24276 51342 24278
rect 51390 24330 51446 24332
rect 51390 24278 51392 24330
rect 51392 24278 51444 24330
rect 51444 24278 51446 24330
rect 51390 24276 51446 24278
rect 51494 24330 51550 24332
rect 51494 24278 51496 24330
rect 51496 24278 51548 24330
rect 51548 24278 51550 24330
rect 51494 24276 51550 24278
rect 50428 22652 50484 22708
rect 51324 23826 51380 23828
rect 51324 23774 51326 23826
rect 51326 23774 51378 23826
rect 51378 23774 51380 23826
rect 51324 23772 51380 23774
rect 51286 22762 51342 22764
rect 51286 22710 51288 22762
rect 51288 22710 51340 22762
rect 51340 22710 51342 22762
rect 51286 22708 51342 22710
rect 51390 22762 51446 22764
rect 51390 22710 51392 22762
rect 51392 22710 51444 22762
rect 51444 22710 51446 22762
rect 51390 22708 51446 22710
rect 51494 22762 51550 22764
rect 51494 22710 51496 22762
rect 51496 22710 51548 22762
rect 51548 22710 51550 22762
rect 51494 22708 51550 22710
rect 51212 21756 51268 21812
rect 51884 23772 51940 23828
rect 52220 23660 52276 23716
rect 52108 23266 52164 23268
rect 52108 23214 52110 23266
rect 52110 23214 52162 23266
rect 52162 23214 52164 23266
rect 52108 23212 52164 23214
rect 50652 20860 50708 20916
rect 50540 18956 50596 19012
rect 50428 16716 50484 16772
rect 50428 15484 50484 15540
rect 50092 15036 50148 15092
rect 50428 15148 50484 15204
rect 49420 14028 49476 14084
rect 49084 13692 49140 13748
rect 44716 11788 44772 11844
rect 45500 12012 45556 12068
rect 43932 11228 43988 11284
rect 44268 11282 44324 11284
rect 44268 11230 44270 11282
rect 44270 11230 44322 11282
rect 44322 11230 44324 11282
rect 44268 11228 44324 11230
rect 45052 11228 45108 11284
rect 43596 11116 43652 11172
rect 43036 10610 43092 10612
rect 43036 10558 43038 10610
rect 43038 10558 43090 10610
rect 43090 10558 43092 10610
rect 43036 10556 43092 10558
rect 42364 9714 42420 9716
rect 42364 9662 42366 9714
rect 42366 9662 42418 9714
rect 42418 9662 42420 9714
rect 42364 9660 42420 9662
rect 42588 9154 42644 9156
rect 42588 9102 42590 9154
rect 42590 9102 42642 9154
rect 42642 9102 42644 9154
rect 42588 9100 42644 9102
rect 42252 8316 42308 8372
rect 42476 8258 42532 8260
rect 42476 8206 42478 8258
rect 42478 8206 42530 8258
rect 42530 8206 42532 8258
rect 42476 8204 42532 8206
rect 42812 9212 42868 9268
rect 42812 8988 42868 9044
rect 41244 7586 41300 7588
rect 41244 7534 41246 7586
rect 41246 7534 41298 7586
rect 41298 7534 41300 7586
rect 41244 7532 41300 7534
rect 42140 7586 42196 7588
rect 42140 7534 42142 7586
rect 42142 7534 42194 7586
rect 42194 7534 42196 7586
rect 42140 7532 42196 7534
rect 41132 7420 41188 7476
rect 42028 7474 42084 7476
rect 42028 7422 42030 7474
rect 42030 7422 42082 7474
rect 42082 7422 42084 7474
rect 42028 7420 42084 7422
rect 40236 6188 40292 6244
rect 39452 5122 39508 5124
rect 39452 5070 39454 5122
rect 39454 5070 39506 5122
rect 39506 5070 39508 5122
rect 39452 5068 39508 5070
rect 42028 6690 42084 6692
rect 42028 6638 42030 6690
rect 42030 6638 42082 6690
rect 42082 6638 42084 6690
rect 42028 6636 42084 6638
rect 42252 6636 42308 6692
rect 43036 9042 43092 9044
rect 43036 8990 43038 9042
rect 43038 8990 43090 9042
rect 43090 8990 43092 9042
rect 43036 8988 43092 8990
rect 43372 9884 43428 9940
rect 43484 9772 43540 9828
rect 44132 11002 44188 11004
rect 44132 10950 44134 11002
rect 44134 10950 44186 11002
rect 44186 10950 44188 11002
rect 44132 10948 44188 10950
rect 44236 11002 44292 11004
rect 44236 10950 44238 11002
rect 44238 10950 44290 11002
rect 44290 10950 44292 11002
rect 44236 10948 44292 10950
rect 44340 11002 44396 11004
rect 44340 10950 44342 11002
rect 44342 10950 44394 11002
rect 44394 10950 44396 11002
rect 44340 10948 44396 10950
rect 45276 11116 45332 11172
rect 45164 9884 45220 9940
rect 43484 9324 43540 9380
rect 44132 9434 44188 9436
rect 44132 9382 44134 9434
rect 44134 9382 44186 9434
rect 44186 9382 44188 9434
rect 44132 9380 44188 9382
rect 44236 9434 44292 9436
rect 44236 9382 44238 9434
rect 44238 9382 44290 9434
rect 44290 9382 44292 9434
rect 44236 9380 44292 9382
rect 44340 9434 44396 9436
rect 44340 9382 44342 9434
rect 44342 9382 44394 9434
rect 44394 9382 44396 9434
rect 44340 9380 44396 9382
rect 45276 9660 45332 9716
rect 44716 9212 44772 9268
rect 45388 9324 45444 9380
rect 44604 8876 44660 8932
rect 43484 8258 43540 8260
rect 43484 8206 43486 8258
rect 43486 8206 43538 8258
rect 43538 8206 43540 8258
rect 43484 8204 43540 8206
rect 43260 7532 43316 7588
rect 43148 6914 43204 6916
rect 43148 6862 43150 6914
rect 43150 6862 43202 6914
rect 43202 6862 43204 6914
rect 43148 6860 43204 6862
rect 43036 6636 43092 6692
rect 41244 5852 41300 5908
rect 40348 5404 40404 5460
rect 40012 5068 40068 5124
rect 40684 5122 40740 5124
rect 40684 5070 40686 5122
rect 40686 5070 40738 5122
rect 40738 5070 40740 5122
rect 40684 5068 40740 5070
rect 40348 4396 40404 4452
rect 41580 5234 41636 5236
rect 41580 5182 41582 5234
rect 41582 5182 41634 5234
rect 41634 5182 41636 5234
rect 41580 5180 41636 5182
rect 41916 4844 41972 4900
rect 38108 3500 38164 3556
rect 41356 4450 41412 4452
rect 41356 4398 41358 4450
rect 41358 4398 41410 4450
rect 41410 4398 41412 4450
rect 41356 4396 41412 4398
rect 41580 4338 41636 4340
rect 41580 4286 41582 4338
rect 41582 4286 41634 4338
rect 41634 4286 41636 4338
rect 41580 4284 41636 4286
rect 41356 3612 41412 3668
rect 41132 3500 41188 3556
rect 41468 3554 41524 3556
rect 41468 3502 41470 3554
rect 41470 3502 41522 3554
rect 41522 3502 41524 3554
rect 41468 3500 41524 3502
rect 42140 5068 42196 5124
rect 42364 3612 42420 3668
rect 43036 6076 43092 6132
rect 42812 5906 42868 5908
rect 42812 5854 42814 5906
rect 42814 5854 42866 5906
rect 42866 5854 42868 5906
rect 42812 5852 42868 5854
rect 44132 7866 44188 7868
rect 44132 7814 44134 7866
rect 44134 7814 44186 7866
rect 44186 7814 44188 7866
rect 44132 7812 44188 7814
rect 44236 7866 44292 7868
rect 44236 7814 44238 7866
rect 44238 7814 44290 7866
rect 44290 7814 44292 7866
rect 44236 7812 44292 7814
rect 44340 7866 44396 7868
rect 44340 7814 44342 7866
rect 44342 7814 44394 7866
rect 44394 7814 44396 7866
rect 44340 7812 44396 7814
rect 44268 7420 44324 7476
rect 43932 6914 43988 6916
rect 43932 6862 43934 6914
rect 43934 6862 43986 6914
rect 43986 6862 43988 6914
rect 43932 6860 43988 6862
rect 45276 9100 45332 9156
rect 45948 11506 46004 11508
rect 45948 11454 45950 11506
rect 45950 11454 46002 11506
rect 46002 11454 46004 11506
rect 45948 11452 46004 11454
rect 46396 10722 46452 10724
rect 46396 10670 46398 10722
rect 46398 10670 46450 10722
rect 46450 10670 46452 10722
rect 46396 10668 46452 10670
rect 47516 11676 47572 11732
rect 46284 10444 46340 10500
rect 46620 10444 46676 10500
rect 47068 11228 47124 11284
rect 48524 12460 48580 12516
rect 48300 12236 48356 12292
rect 48300 11900 48356 11956
rect 48076 11228 48132 11284
rect 47964 11116 48020 11172
rect 47852 10668 47908 10724
rect 47068 10444 47124 10500
rect 46956 9938 47012 9940
rect 46956 9886 46958 9938
rect 46958 9886 47010 9938
rect 47010 9886 47012 9938
rect 46956 9884 47012 9886
rect 46508 9714 46564 9716
rect 46508 9662 46510 9714
rect 46510 9662 46562 9714
rect 46562 9662 46564 9714
rect 46508 9660 46564 9662
rect 47404 10444 47460 10500
rect 46732 9100 46788 9156
rect 47964 10050 48020 10052
rect 47964 9998 47966 10050
rect 47966 9998 48018 10050
rect 48018 9998 48020 10050
rect 47964 9996 48020 9998
rect 47628 9772 47684 9828
rect 47628 9548 47684 9604
rect 48636 12124 48692 12180
rect 49420 13468 49476 13524
rect 49868 14028 49924 14084
rect 50428 14700 50484 14756
rect 51286 21194 51342 21196
rect 51286 21142 51288 21194
rect 51288 21142 51340 21194
rect 51340 21142 51342 21194
rect 51286 21140 51342 21142
rect 51390 21194 51446 21196
rect 51390 21142 51392 21194
rect 51392 21142 51444 21194
rect 51444 21142 51446 21194
rect 51390 21140 51446 21142
rect 51494 21194 51550 21196
rect 51494 21142 51496 21194
rect 51496 21142 51548 21194
rect 51548 21142 51550 21194
rect 51494 21140 51550 21142
rect 50764 20748 50820 20804
rect 50876 20188 50932 20244
rect 51100 19740 51156 19796
rect 51286 19626 51342 19628
rect 51286 19574 51288 19626
rect 51288 19574 51340 19626
rect 51340 19574 51342 19626
rect 51286 19572 51342 19574
rect 51390 19626 51446 19628
rect 51390 19574 51392 19626
rect 51392 19574 51444 19626
rect 51444 19574 51446 19626
rect 51390 19572 51446 19574
rect 51494 19626 51550 19628
rect 51494 19574 51496 19626
rect 51496 19574 51548 19626
rect 51548 19574 51550 19626
rect 51494 19572 51550 19574
rect 51996 21532 52052 21588
rect 51772 19292 51828 19348
rect 51884 20860 51940 20916
rect 50876 19234 50932 19236
rect 50876 19182 50878 19234
rect 50878 19182 50930 19234
rect 50930 19182 50932 19234
rect 50876 19180 50932 19182
rect 52444 23266 52500 23268
rect 52444 23214 52446 23266
rect 52446 23214 52498 23266
rect 52498 23214 52500 23266
rect 52444 23212 52500 23214
rect 53004 25452 53060 25508
rect 52892 23772 52948 23828
rect 52332 22876 52388 22932
rect 52108 20972 52164 21028
rect 52220 20690 52276 20692
rect 52220 20638 52222 20690
rect 52222 20638 52274 20690
rect 52274 20638 52276 20690
rect 52220 20636 52276 20638
rect 51286 18058 51342 18060
rect 51286 18006 51288 18058
rect 51288 18006 51340 18058
rect 51340 18006 51342 18058
rect 51286 18004 51342 18006
rect 51390 18058 51446 18060
rect 51390 18006 51392 18058
rect 51392 18006 51444 18058
rect 51444 18006 51446 18058
rect 51390 18004 51446 18006
rect 51494 18058 51550 18060
rect 51494 18006 51496 18058
rect 51496 18006 51548 18058
rect 51548 18006 51550 18058
rect 51494 18004 51550 18006
rect 50652 15820 50708 15876
rect 50988 16994 51044 16996
rect 50988 16942 50990 16994
rect 50990 16942 51042 16994
rect 51042 16942 51044 16994
rect 50988 16940 51044 16942
rect 51660 17442 51716 17444
rect 51660 17390 51662 17442
rect 51662 17390 51714 17442
rect 51714 17390 51716 17442
rect 51660 17388 51716 17390
rect 51548 16716 51604 16772
rect 51286 16490 51342 16492
rect 51286 16438 51288 16490
rect 51288 16438 51340 16490
rect 51340 16438 51342 16490
rect 51286 16436 51342 16438
rect 51390 16490 51446 16492
rect 51390 16438 51392 16490
rect 51392 16438 51444 16490
rect 51444 16438 51446 16490
rect 51390 16436 51446 16438
rect 51494 16490 51550 16492
rect 51494 16438 51496 16490
rect 51496 16438 51548 16490
rect 51548 16438 51550 16490
rect 51494 16436 51550 16438
rect 53676 25452 53732 25508
rect 56588 25564 56644 25620
rect 55468 25506 55524 25508
rect 55468 25454 55470 25506
rect 55470 25454 55522 25506
rect 55522 25454 55524 25506
rect 55468 25452 55524 25454
rect 58439 25114 58495 25116
rect 58439 25062 58441 25114
rect 58441 25062 58493 25114
rect 58493 25062 58495 25114
rect 58439 25060 58495 25062
rect 58543 25114 58599 25116
rect 58543 25062 58545 25114
rect 58545 25062 58597 25114
rect 58597 25062 58599 25114
rect 58543 25060 58599 25062
rect 58647 25114 58703 25116
rect 58647 25062 58649 25114
rect 58649 25062 58701 25114
rect 58701 25062 58703 25114
rect 58647 25060 58703 25062
rect 54908 23884 54964 23940
rect 53564 23660 53620 23716
rect 52668 23378 52724 23380
rect 52668 23326 52670 23378
rect 52670 23326 52722 23378
rect 52722 23326 52724 23378
rect 52668 23324 52724 23326
rect 53228 23212 53284 23268
rect 53004 22876 53060 22932
rect 52780 22540 52836 22596
rect 53004 22428 53060 22484
rect 52892 22146 52948 22148
rect 52892 22094 52894 22146
rect 52894 22094 52946 22146
rect 52946 22094 52948 22146
rect 52892 22092 52948 22094
rect 52668 20412 52724 20468
rect 53340 22316 53396 22372
rect 54572 23548 54628 23604
rect 53452 22204 53508 22260
rect 52780 19964 52836 20020
rect 52892 20188 52948 20244
rect 52444 19740 52500 19796
rect 52332 18562 52388 18564
rect 52332 18510 52334 18562
rect 52334 18510 52386 18562
rect 52386 18510 52388 18562
rect 52332 18508 52388 18510
rect 52556 18450 52612 18452
rect 52556 18398 52558 18450
rect 52558 18398 52610 18450
rect 52610 18398 52612 18450
rect 52556 18396 52612 18398
rect 53228 20578 53284 20580
rect 53228 20526 53230 20578
rect 53230 20526 53282 20578
rect 53282 20526 53284 20578
rect 53228 20524 53284 20526
rect 53788 22316 53844 22372
rect 53564 21644 53620 21700
rect 53676 22258 53732 22260
rect 53676 22206 53678 22258
rect 53678 22206 53730 22258
rect 53730 22206 53732 22258
rect 53676 22204 53732 22206
rect 54348 22204 54404 22260
rect 54124 21756 54180 21812
rect 53900 21532 53956 21588
rect 53340 20188 53396 20244
rect 53452 20748 53508 20804
rect 54012 20130 54068 20132
rect 54012 20078 54014 20130
rect 54014 20078 54066 20130
rect 54066 20078 54068 20130
rect 54012 20076 54068 20078
rect 53004 19180 53060 19236
rect 53340 19292 53396 19348
rect 53228 17836 53284 17892
rect 51996 17388 52052 17444
rect 51772 16716 51828 16772
rect 51436 16210 51492 16212
rect 51436 16158 51438 16210
rect 51438 16158 51490 16210
rect 51490 16158 51492 16210
rect 51436 16156 51492 16158
rect 51436 15372 51492 15428
rect 50652 15260 50708 15316
rect 51212 15314 51268 15316
rect 51212 15262 51214 15314
rect 51214 15262 51266 15314
rect 51266 15262 51268 15314
rect 51212 15260 51268 15262
rect 51660 16044 51716 16100
rect 51884 16044 51940 16100
rect 52108 16940 52164 16996
rect 51772 15932 51828 15988
rect 53116 17778 53172 17780
rect 53116 17726 53118 17778
rect 53118 17726 53170 17778
rect 53170 17726 53172 17778
rect 53116 17724 53172 17726
rect 54460 19292 54516 19348
rect 53900 18284 53956 18340
rect 54460 18562 54516 18564
rect 54460 18510 54462 18562
rect 54462 18510 54514 18562
rect 54514 18510 54516 18562
rect 54460 18508 54516 18510
rect 54796 21532 54852 21588
rect 55132 22316 55188 22372
rect 54796 20914 54852 20916
rect 54796 20862 54798 20914
rect 54798 20862 54850 20914
rect 54850 20862 54852 20914
rect 54796 20860 54852 20862
rect 55020 20802 55076 20804
rect 55020 20750 55022 20802
rect 55022 20750 55074 20802
rect 55074 20750 55076 20802
rect 55020 20748 55076 20750
rect 55580 23938 55636 23940
rect 55580 23886 55582 23938
rect 55582 23886 55634 23938
rect 55634 23886 55636 23938
rect 55580 23884 55636 23886
rect 55804 23324 55860 23380
rect 55468 23266 55524 23268
rect 55468 23214 55470 23266
rect 55470 23214 55522 23266
rect 55522 23214 55524 23266
rect 55468 23212 55524 23214
rect 55356 21756 55412 21812
rect 55244 21586 55300 21588
rect 55244 21534 55246 21586
rect 55246 21534 55298 21586
rect 55298 21534 55300 21586
rect 55244 21532 55300 21534
rect 55468 21644 55524 21700
rect 56364 22370 56420 22372
rect 56364 22318 56366 22370
rect 56366 22318 56418 22370
rect 56418 22318 56420 22370
rect 56364 22316 56420 22318
rect 55804 21586 55860 21588
rect 55804 21534 55806 21586
rect 55806 21534 55858 21586
rect 55858 21534 55860 21586
rect 55804 21532 55860 21534
rect 55244 20076 55300 20132
rect 54796 19180 54852 19236
rect 54908 18732 54964 18788
rect 54236 18284 54292 18340
rect 53564 17724 53620 17780
rect 53564 17052 53620 17108
rect 53340 16716 53396 16772
rect 53228 16156 53284 16212
rect 51772 15260 51828 15316
rect 53452 15314 53508 15316
rect 53452 15262 53454 15314
rect 53454 15262 53506 15314
rect 53506 15262 53508 15314
rect 53452 15260 53508 15262
rect 51286 14922 51342 14924
rect 51286 14870 51288 14922
rect 51288 14870 51340 14922
rect 51340 14870 51342 14922
rect 51286 14868 51342 14870
rect 51390 14922 51446 14924
rect 51390 14870 51392 14922
rect 51392 14870 51444 14922
rect 51444 14870 51446 14922
rect 51390 14868 51446 14870
rect 51494 14922 51550 14924
rect 51494 14870 51496 14922
rect 51496 14870 51548 14922
rect 51548 14870 51550 14922
rect 51494 14868 51550 14870
rect 50316 13692 50372 13748
rect 49420 12178 49476 12180
rect 49420 12126 49422 12178
rect 49422 12126 49474 12178
rect 49474 12126 49476 12178
rect 49420 12124 49476 12126
rect 48860 10722 48916 10724
rect 48860 10670 48862 10722
rect 48862 10670 48914 10722
rect 48914 10670 48916 10722
rect 48860 10668 48916 10670
rect 48636 10444 48692 10500
rect 45500 8764 45556 8820
rect 45948 8764 46004 8820
rect 45388 8204 45444 8260
rect 45276 7980 45332 8036
rect 45052 7586 45108 7588
rect 45052 7534 45054 7586
rect 45054 7534 45106 7586
rect 45106 7534 45108 7586
rect 45052 7532 45108 7534
rect 46732 8034 46788 8036
rect 46732 7982 46734 8034
rect 46734 7982 46786 8034
rect 46786 7982 46788 8034
rect 46732 7980 46788 7982
rect 43708 6748 43764 6804
rect 44268 6690 44324 6692
rect 44268 6638 44270 6690
rect 44270 6638 44322 6690
rect 44322 6638 44324 6690
rect 44268 6636 44324 6638
rect 43596 6412 43652 6468
rect 44132 6298 44188 6300
rect 44132 6246 44134 6298
rect 44134 6246 44186 6298
rect 44186 6246 44188 6298
rect 44132 6244 44188 6246
rect 44236 6298 44292 6300
rect 44236 6246 44238 6298
rect 44238 6246 44290 6298
rect 44290 6246 44292 6298
rect 44236 6244 44292 6246
rect 44340 6298 44396 6300
rect 44340 6246 44342 6298
rect 44342 6246 44394 6298
rect 44394 6246 44396 6298
rect 44340 6244 44396 6246
rect 43820 5122 43876 5124
rect 43820 5070 43822 5122
rect 43822 5070 43874 5122
rect 43874 5070 43876 5122
rect 43820 5068 43876 5070
rect 44132 4730 44188 4732
rect 44132 4678 44134 4730
rect 44134 4678 44186 4730
rect 44186 4678 44188 4730
rect 44132 4676 44188 4678
rect 44236 4730 44292 4732
rect 44236 4678 44238 4730
rect 44238 4678 44290 4730
rect 44290 4678 44292 4730
rect 44236 4676 44292 4678
rect 44340 4730 44396 4732
rect 44340 4678 44342 4730
rect 44342 4678 44394 4730
rect 44394 4678 44396 4730
rect 44340 4676 44396 4678
rect 43708 4620 43764 4676
rect 43932 4396 43988 4452
rect 44156 4338 44212 4340
rect 44156 4286 44158 4338
rect 44158 4286 44210 4338
rect 44210 4286 44212 4338
rect 44156 4284 44212 4286
rect 44828 6860 44884 6916
rect 45388 6748 45444 6804
rect 44828 5852 44884 5908
rect 45724 6524 45780 6580
rect 45388 5740 45444 5796
rect 46284 7474 46340 7476
rect 46284 7422 46286 7474
rect 46286 7422 46338 7474
rect 46338 7422 46340 7474
rect 46284 7420 46340 7422
rect 46060 6690 46116 6692
rect 46060 6638 46062 6690
rect 46062 6638 46114 6690
rect 46114 6638 46116 6690
rect 46060 6636 46116 6638
rect 46508 6524 46564 6580
rect 45836 6412 45892 6468
rect 46844 6636 46900 6692
rect 46732 6412 46788 6468
rect 47516 8818 47572 8820
rect 47516 8766 47518 8818
rect 47518 8766 47570 8818
rect 47570 8766 47572 8818
rect 47516 8764 47572 8766
rect 48412 9548 48468 9604
rect 48188 9042 48244 9044
rect 48188 8990 48190 9042
rect 48190 8990 48242 9042
rect 48242 8990 48244 9042
rect 48188 8988 48244 8990
rect 48412 8258 48468 8260
rect 48412 8206 48414 8258
rect 48414 8206 48466 8258
rect 48466 8206 48468 8258
rect 48412 8204 48468 8206
rect 48076 7980 48132 8036
rect 47180 6524 47236 6580
rect 45836 5180 45892 5236
rect 47740 6300 47796 6356
rect 45612 5122 45668 5124
rect 45612 5070 45614 5122
rect 45614 5070 45666 5122
rect 45666 5070 45668 5122
rect 45612 5068 45668 5070
rect 44940 4732 44996 4788
rect 46844 5068 46900 5124
rect 46732 4732 46788 4788
rect 45164 4450 45220 4452
rect 45164 4398 45166 4450
rect 45166 4398 45218 4450
rect 45218 4398 45220 4450
rect 45164 4396 45220 4398
rect 46732 4396 46788 4452
rect 47404 4450 47460 4452
rect 47404 4398 47406 4450
rect 47406 4398 47458 4450
rect 47458 4398 47460 4450
rect 47404 4396 47460 4398
rect 48300 6636 48356 6692
rect 48076 6018 48132 6020
rect 48076 5966 48078 6018
rect 48078 5966 48130 6018
rect 48130 5966 48132 6018
rect 48076 5964 48132 5966
rect 48076 5292 48132 5348
rect 49084 11954 49140 11956
rect 49084 11902 49086 11954
rect 49086 11902 49138 11954
rect 49138 11902 49140 11954
rect 49084 11900 49140 11902
rect 49084 11676 49140 11732
rect 49644 12348 49700 12404
rect 50204 13132 50260 13188
rect 50092 12402 50148 12404
rect 50092 12350 50094 12402
rect 50094 12350 50146 12402
rect 50146 12350 50148 12402
rect 50092 12348 50148 12350
rect 49868 11676 49924 11732
rect 49980 12124 50036 12180
rect 49644 11004 49700 11060
rect 50316 11506 50372 11508
rect 50316 11454 50318 11506
rect 50318 11454 50370 11506
rect 50370 11454 50372 11506
rect 50316 11452 50372 11454
rect 50540 14306 50596 14308
rect 50540 14254 50542 14306
rect 50542 14254 50594 14306
rect 50594 14254 50596 14306
rect 50540 14252 50596 14254
rect 51100 13804 51156 13860
rect 50988 12908 51044 12964
rect 51212 13468 51268 13524
rect 51286 13354 51342 13356
rect 51286 13302 51288 13354
rect 51288 13302 51340 13354
rect 51340 13302 51342 13354
rect 51286 13300 51342 13302
rect 51390 13354 51446 13356
rect 51390 13302 51392 13354
rect 51392 13302 51444 13354
rect 51444 13302 51446 13354
rect 51390 13300 51446 13302
rect 51494 13354 51550 13356
rect 51494 13302 51496 13354
rect 51496 13302 51548 13354
rect 51548 13302 51550 13354
rect 51494 13300 51550 13302
rect 51660 13132 51716 13188
rect 51436 13074 51492 13076
rect 51436 13022 51438 13074
rect 51438 13022 51490 13074
rect 51490 13022 51492 13074
rect 51436 13020 51492 13022
rect 51324 12962 51380 12964
rect 51324 12910 51326 12962
rect 51326 12910 51378 12962
rect 51378 12910 51380 12962
rect 51324 12908 51380 12910
rect 51548 12850 51604 12852
rect 51548 12798 51550 12850
rect 51550 12798 51602 12850
rect 51602 12798 51604 12850
rect 51548 12796 51604 12798
rect 51660 12290 51716 12292
rect 51660 12238 51662 12290
rect 51662 12238 51714 12290
rect 51714 12238 51716 12290
rect 51660 12236 51716 12238
rect 51100 12178 51156 12180
rect 51100 12126 51102 12178
rect 51102 12126 51154 12178
rect 51154 12126 51156 12178
rect 51100 12124 51156 12126
rect 51548 12066 51604 12068
rect 51548 12014 51550 12066
rect 51550 12014 51602 12066
rect 51602 12014 51604 12066
rect 51548 12012 51604 12014
rect 51286 11786 51342 11788
rect 51286 11734 51288 11786
rect 51288 11734 51340 11786
rect 51340 11734 51342 11786
rect 51286 11732 51342 11734
rect 51390 11786 51446 11788
rect 51390 11734 51392 11786
rect 51392 11734 51444 11786
rect 51444 11734 51446 11786
rect 51390 11732 51446 11734
rect 51494 11786 51550 11788
rect 51494 11734 51496 11786
rect 51496 11734 51548 11786
rect 51548 11734 51550 11786
rect 51494 11732 51550 11734
rect 50764 11564 50820 11620
rect 53452 14812 53508 14868
rect 51772 11506 51828 11508
rect 51772 11454 51774 11506
rect 51774 11454 51826 11506
rect 51826 11454 51828 11506
rect 51772 11452 51828 11454
rect 51884 14700 51940 14756
rect 50652 11004 50708 11060
rect 49644 10556 49700 10612
rect 49308 10220 49364 10276
rect 50428 10498 50484 10500
rect 50428 10446 50430 10498
rect 50430 10446 50482 10498
rect 50482 10446 50484 10498
rect 50428 10444 50484 10446
rect 49980 9996 50036 10052
rect 49532 9772 49588 9828
rect 49868 9660 49924 9716
rect 48748 8876 48804 8932
rect 48972 8988 49028 9044
rect 48748 8258 48804 8260
rect 48748 8206 48750 8258
rect 48750 8206 48802 8258
rect 48802 8206 48804 8258
rect 48748 8204 48804 8206
rect 48972 6690 49028 6692
rect 48972 6638 48974 6690
rect 48974 6638 49026 6690
rect 49026 6638 49028 6690
rect 48972 6636 49028 6638
rect 48860 6524 48916 6580
rect 48748 6300 48804 6356
rect 48972 5906 49028 5908
rect 48972 5854 48974 5906
rect 48974 5854 49026 5906
rect 49026 5854 49028 5906
rect 48972 5852 49028 5854
rect 48860 5292 48916 5348
rect 49084 5404 49140 5460
rect 48076 4226 48132 4228
rect 48076 4174 48078 4226
rect 48078 4174 48130 4226
rect 48130 4174 48132 4226
rect 48076 4172 48132 4174
rect 49196 5346 49252 5348
rect 49196 5294 49198 5346
rect 49198 5294 49250 5346
rect 49250 5294 49252 5346
rect 49196 5292 49252 5294
rect 49532 6524 49588 6580
rect 50652 10444 50708 10500
rect 51286 10218 51342 10220
rect 51286 10166 51288 10218
rect 51288 10166 51340 10218
rect 51340 10166 51342 10218
rect 51286 10164 51342 10166
rect 51390 10218 51446 10220
rect 51390 10166 51392 10218
rect 51392 10166 51444 10218
rect 51444 10166 51446 10218
rect 51390 10164 51446 10166
rect 51494 10218 51550 10220
rect 51494 10166 51496 10218
rect 51496 10166 51548 10218
rect 51548 10166 51550 10218
rect 51494 10164 51550 10166
rect 51660 9884 51716 9940
rect 49980 8876 50036 8932
rect 50764 9042 50820 9044
rect 50764 8990 50766 9042
rect 50766 8990 50818 9042
rect 50818 8990 50820 9042
rect 50764 8988 50820 8990
rect 51324 8930 51380 8932
rect 51324 8878 51326 8930
rect 51326 8878 51378 8930
rect 51378 8878 51380 8930
rect 51324 8876 51380 8878
rect 51772 8876 51828 8932
rect 51286 8650 51342 8652
rect 51286 8598 51288 8650
rect 51288 8598 51340 8650
rect 51340 8598 51342 8650
rect 51286 8596 51342 8598
rect 51390 8650 51446 8652
rect 51390 8598 51392 8650
rect 51392 8598 51444 8650
rect 51444 8598 51446 8650
rect 51390 8596 51446 8598
rect 51494 8650 51550 8652
rect 51494 8598 51496 8650
rect 51496 8598 51548 8650
rect 51548 8598 51550 8650
rect 51494 8596 51550 8598
rect 51286 7082 51342 7084
rect 51286 7030 51288 7082
rect 51288 7030 51340 7082
rect 51340 7030 51342 7082
rect 51286 7028 51342 7030
rect 51390 7082 51446 7084
rect 51390 7030 51392 7082
rect 51392 7030 51444 7082
rect 51444 7030 51446 7082
rect 51390 7028 51446 7030
rect 51494 7082 51550 7084
rect 51494 7030 51496 7082
rect 51496 7030 51548 7082
rect 51548 7030 51550 7082
rect 51494 7028 51550 7030
rect 50092 6018 50148 6020
rect 50092 5966 50094 6018
rect 50094 5966 50146 6018
rect 50146 5966 50148 6018
rect 50092 5964 50148 5966
rect 50316 6188 50372 6244
rect 51100 6636 51156 6692
rect 51548 6636 51604 6692
rect 51324 6524 51380 6580
rect 50764 6076 50820 6132
rect 50988 6188 51044 6244
rect 52108 14306 52164 14308
rect 52108 14254 52110 14306
rect 52110 14254 52162 14306
rect 52162 14254 52164 14306
rect 52108 14252 52164 14254
rect 52556 12908 52612 12964
rect 51996 12850 52052 12852
rect 51996 12798 51998 12850
rect 51998 12798 52050 12850
rect 52050 12798 52052 12850
rect 51996 12796 52052 12798
rect 52668 13132 52724 13188
rect 53004 14252 53060 14308
rect 53228 14028 53284 14084
rect 53116 13468 53172 13524
rect 53676 16156 53732 16212
rect 54012 17836 54068 17892
rect 53900 16994 53956 16996
rect 53900 16942 53902 16994
rect 53902 16942 53954 16994
rect 53954 16942 53956 16994
rect 53900 16940 53956 16942
rect 53788 15148 53844 15204
rect 53900 16716 53956 16772
rect 54236 17388 54292 17444
rect 54572 17836 54628 17892
rect 55132 18508 55188 18564
rect 54796 17276 54852 17332
rect 54348 16044 54404 16100
rect 54012 15148 54068 15204
rect 53900 14924 53956 14980
rect 53564 13020 53620 13076
rect 53788 14252 53844 14308
rect 53788 13020 53844 13076
rect 52108 12290 52164 12292
rect 52108 12238 52110 12290
rect 52110 12238 52162 12290
rect 52162 12238 52164 12290
rect 52108 12236 52164 12238
rect 53676 12962 53732 12964
rect 53676 12910 53678 12962
rect 53678 12910 53730 12962
rect 53730 12910 53732 12962
rect 53676 12908 53732 12910
rect 53228 12796 53284 12852
rect 53340 12684 53396 12740
rect 53116 11564 53172 11620
rect 53228 11676 53284 11732
rect 53228 11340 53284 11396
rect 52108 8316 52164 8372
rect 52892 8204 52948 8260
rect 53004 8316 53060 8372
rect 52780 6914 52836 6916
rect 52780 6862 52782 6914
rect 52782 6862 52834 6914
rect 52834 6862 52836 6914
rect 52780 6860 52836 6862
rect 53788 11900 53844 11956
rect 54572 16268 54628 16324
rect 54684 16156 54740 16212
rect 55020 16380 55076 16436
rect 55244 17388 55300 17444
rect 55356 17276 55412 17332
rect 55692 20636 55748 20692
rect 56028 21420 56084 21476
rect 56700 21474 56756 21476
rect 56700 21422 56702 21474
rect 56702 21422 56754 21474
rect 56754 21422 56756 21474
rect 56700 21420 56756 21422
rect 56140 20636 56196 20692
rect 55580 16716 55636 16772
rect 54908 16098 54964 16100
rect 54908 16046 54910 16098
rect 54910 16046 54962 16098
rect 54962 16046 54964 16098
rect 54908 16044 54964 16046
rect 55356 16044 55412 16100
rect 55020 15986 55076 15988
rect 55020 15934 55022 15986
rect 55022 15934 55074 15986
rect 55074 15934 55076 15986
rect 55020 15932 55076 15934
rect 54796 15484 54852 15540
rect 55468 16380 55524 16436
rect 55244 15538 55300 15540
rect 55244 15486 55246 15538
rect 55246 15486 55298 15538
rect 55298 15486 55300 15538
rect 55244 15484 55300 15486
rect 55132 15260 55188 15316
rect 54572 14924 54628 14980
rect 54572 14306 54628 14308
rect 54572 14254 54574 14306
rect 54574 14254 54626 14306
rect 54626 14254 54628 14306
rect 54572 14252 54628 14254
rect 54684 13692 54740 13748
rect 55132 14812 55188 14868
rect 55692 16268 55748 16324
rect 55580 16210 55636 16212
rect 55580 16158 55582 16210
rect 55582 16158 55634 16210
rect 55634 16158 55636 16210
rect 55580 16156 55636 16158
rect 56924 23212 56980 23268
rect 57036 23324 57092 23380
rect 57708 23884 57764 23940
rect 57596 23714 57652 23716
rect 57596 23662 57598 23714
rect 57598 23662 57650 23714
rect 57650 23662 57652 23714
rect 57596 23660 57652 23662
rect 57932 23548 57988 23604
rect 58439 23546 58495 23548
rect 58439 23494 58441 23546
rect 58441 23494 58493 23546
rect 58493 23494 58495 23546
rect 58439 23492 58495 23494
rect 58543 23546 58599 23548
rect 58543 23494 58545 23546
rect 58545 23494 58597 23546
rect 58597 23494 58599 23546
rect 58543 23492 58599 23494
rect 58647 23546 58703 23548
rect 58647 23494 58649 23546
rect 58649 23494 58701 23546
rect 58701 23494 58703 23546
rect 58647 23492 58703 23494
rect 58439 21978 58495 21980
rect 58439 21926 58441 21978
rect 58441 21926 58493 21978
rect 58493 21926 58495 21978
rect 58439 21924 58495 21926
rect 58543 21978 58599 21980
rect 58543 21926 58545 21978
rect 58545 21926 58597 21978
rect 58597 21926 58599 21978
rect 58543 21924 58599 21926
rect 58647 21978 58703 21980
rect 58647 21926 58649 21978
rect 58649 21926 58701 21978
rect 58701 21926 58703 21978
rect 58647 21924 58703 21926
rect 57932 21586 57988 21588
rect 57932 21534 57934 21586
rect 57934 21534 57986 21586
rect 57986 21534 57988 21586
rect 57932 21532 57988 21534
rect 55356 14364 55412 14420
rect 55244 14028 55300 14084
rect 54908 13132 54964 13188
rect 54460 12962 54516 12964
rect 54460 12910 54462 12962
rect 54462 12910 54514 12962
rect 54514 12910 54516 12962
rect 54460 12908 54516 12910
rect 54012 12738 54068 12740
rect 54012 12686 54014 12738
rect 54014 12686 54066 12738
rect 54066 12686 54068 12738
rect 54012 12684 54068 12686
rect 55132 12908 55188 12964
rect 55356 13746 55412 13748
rect 55356 13694 55358 13746
rect 55358 13694 55410 13746
rect 55410 13694 55412 13746
rect 55356 13692 55412 13694
rect 55468 13074 55524 13076
rect 55468 13022 55470 13074
rect 55470 13022 55522 13074
rect 55522 13022 55524 13074
rect 55468 13020 55524 13022
rect 55468 12684 55524 12740
rect 54908 12348 54964 12404
rect 53900 11676 53956 11732
rect 53564 11564 53620 11620
rect 54236 11452 54292 11508
rect 55356 12402 55412 12404
rect 55356 12350 55358 12402
rect 55358 12350 55410 12402
rect 55410 12350 55412 12402
rect 55356 12348 55412 12350
rect 54796 12178 54852 12180
rect 54796 12126 54798 12178
rect 54798 12126 54850 12178
rect 54850 12126 54852 12178
rect 54796 12124 54852 12126
rect 55804 14476 55860 14532
rect 56252 14812 56308 14868
rect 56140 14028 56196 14084
rect 55916 13970 55972 13972
rect 55916 13918 55918 13970
rect 55918 13918 55970 13970
rect 55970 13918 55972 13970
rect 55916 13916 55972 13918
rect 55692 13692 55748 13748
rect 55692 13132 55748 13188
rect 57708 20130 57764 20132
rect 57708 20078 57710 20130
rect 57710 20078 57762 20130
rect 57762 20078 57764 20130
rect 57708 20076 57764 20078
rect 58439 20410 58495 20412
rect 58439 20358 58441 20410
rect 58441 20358 58493 20410
rect 58493 20358 58495 20410
rect 58439 20356 58495 20358
rect 58543 20410 58599 20412
rect 58543 20358 58545 20410
rect 58545 20358 58597 20410
rect 58597 20358 58599 20410
rect 58543 20356 58599 20358
rect 58647 20410 58703 20412
rect 58647 20358 58649 20410
rect 58649 20358 58701 20410
rect 58701 20358 58703 20410
rect 58647 20356 58703 20358
rect 58044 19180 58100 19236
rect 57484 18732 57540 18788
rect 58439 18842 58495 18844
rect 58439 18790 58441 18842
rect 58441 18790 58493 18842
rect 58493 18790 58495 18842
rect 58439 18788 58495 18790
rect 58543 18842 58599 18844
rect 58543 18790 58545 18842
rect 58545 18790 58597 18842
rect 58597 18790 58599 18842
rect 58543 18788 58599 18790
rect 58647 18842 58703 18844
rect 58647 18790 58649 18842
rect 58649 18790 58701 18842
rect 58701 18790 58703 18842
rect 58647 18788 58703 18790
rect 57036 17442 57092 17444
rect 57036 17390 57038 17442
rect 57038 17390 57090 17442
rect 57090 17390 57092 17442
rect 57036 17388 57092 17390
rect 56476 16828 56532 16884
rect 58439 17274 58495 17276
rect 58439 17222 58441 17274
rect 58441 17222 58493 17274
rect 58493 17222 58495 17274
rect 58439 17220 58495 17222
rect 58543 17274 58599 17276
rect 58543 17222 58545 17274
rect 58545 17222 58597 17274
rect 58597 17222 58599 17274
rect 58543 17220 58599 17222
rect 58647 17274 58703 17276
rect 58647 17222 58649 17274
rect 58649 17222 58701 17274
rect 58701 17222 58703 17274
rect 58647 17220 58703 17222
rect 58156 17052 58212 17108
rect 56924 16770 56980 16772
rect 56924 16718 56926 16770
rect 56926 16718 56978 16770
rect 56978 16718 56980 16770
rect 56924 16716 56980 16718
rect 57148 16604 57204 16660
rect 56476 14530 56532 14532
rect 56476 14478 56478 14530
rect 56478 14478 56530 14530
rect 56530 14478 56532 14530
rect 56476 14476 56532 14478
rect 55804 13020 55860 13076
rect 56028 13132 56084 13188
rect 56028 12684 56084 12740
rect 55916 12572 55972 12628
rect 55692 12290 55748 12292
rect 55692 12238 55694 12290
rect 55694 12238 55746 12290
rect 55746 12238 55748 12290
rect 55692 12236 55748 12238
rect 55020 11900 55076 11956
rect 55244 11900 55300 11956
rect 55244 11452 55300 11508
rect 55132 11394 55188 11396
rect 55132 11342 55134 11394
rect 55134 11342 55186 11394
rect 55186 11342 55188 11394
rect 55132 11340 55188 11342
rect 54236 10386 54292 10388
rect 54236 10334 54238 10386
rect 54238 10334 54290 10386
rect 54290 10334 54292 10386
rect 54236 10332 54292 10334
rect 54684 9884 54740 9940
rect 54572 9602 54628 9604
rect 54572 9550 54574 9602
rect 54574 9550 54626 9602
rect 54626 9550 54628 9602
rect 54572 9548 54628 9550
rect 54348 9324 54404 9380
rect 54908 9714 54964 9716
rect 54908 9662 54910 9714
rect 54910 9662 54962 9714
rect 54962 9662 54964 9714
rect 54908 9660 54964 9662
rect 54796 8988 54852 9044
rect 53564 8930 53620 8932
rect 53564 8878 53566 8930
rect 53566 8878 53618 8930
rect 53618 8878 53620 8930
rect 53564 8876 53620 8878
rect 53228 6748 53284 6804
rect 52108 6636 52164 6692
rect 51996 6466 52052 6468
rect 51996 6414 51998 6466
rect 51998 6414 52050 6466
rect 52050 6414 52052 6466
rect 51996 6412 52052 6414
rect 51884 6188 51940 6244
rect 51100 6018 51156 6020
rect 51100 5966 51102 6018
rect 51102 5966 51154 6018
rect 51154 5966 51156 6018
rect 51100 5964 51156 5966
rect 52668 6578 52724 6580
rect 52668 6526 52670 6578
rect 52670 6526 52722 6578
rect 52722 6526 52724 6578
rect 52668 6524 52724 6526
rect 52220 6130 52276 6132
rect 52220 6078 52222 6130
rect 52222 6078 52274 6130
rect 52274 6078 52276 6130
rect 52220 6076 52276 6078
rect 52780 6076 52836 6132
rect 53900 6412 53956 6468
rect 54908 8428 54964 8484
rect 54796 8316 54852 8372
rect 55468 11170 55524 11172
rect 55468 11118 55470 11170
rect 55470 11118 55522 11170
rect 55522 11118 55524 11170
rect 55468 11116 55524 11118
rect 55468 10780 55524 10836
rect 55916 11394 55972 11396
rect 55916 11342 55918 11394
rect 55918 11342 55970 11394
rect 55970 11342 55972 11394
rect 55916 11340 55972 11342
rect 57596 16658 57652 16660
rect 57596 16606 57598 16658
rect 57598 16606 57650 16658
rect 57650 16606 57652 16658
rect 57596 16604 57652 16606
rect 57372 16098 57428 16100
rect 57372 16046 57374 16098
rect 57374 16046 57426 16098
rect 57426 16046 57428 16098
rect 57372 16044 57428 16046
rect 57932 16882 57988 16884
rect 57932 16830 57934 16882
rect 57934 16830 57986 16882
rect 57986 16830 57988 16882
rect 57932 16828 57988 16830
rect 58044 16604 58100 16660
rect 58439 15706 58495 15708
rect 58439 15654 58441 15706
rect 58441 15654 58493 15706
rect 58493 15654 58495 15706
rect 58439 15652 58495 15654
rect 58543 15706 58599 15708
rect 58543 15654 58545 15706
rect 58545 15654 58597 15706
rect 58597 15654 58599 15706
rect 58543 15652 58599 15654
rect 58647 15706 58703 15708
rect 58647 15654 58649 15706
rect 58649 15654 58701 15706
rect 58701 15654 58703 15706
rect 58647 15652 58703 15654
rect 57260 14476 57316 14532
rect 57036 14418 57092 14420
rect 57036 14366 57038 14418
rect 57038 14366 57090 14418
rect 57090 14366 57092 14418
rect 57036 14364 57092 14366
rect 57260 13132 57316 13188
rect 56700 13020 56756 13076
rect 56476 12962 56532 12964
rect 56476 12910 56478 12962
rect 56478 12910 56530 12962
rect 56530 12910 56532 12962
rect 56476 12908 56532 12910
rect 56700 12348 56756 12404
rect 56700 11900 56756 11956
rect 57148 12738 57204 12740
rect 57148 12686 57150 12738
rect 57150 12686 57202 12738
rect 57202 12686 57204 12738
rect 57148 12684 57204 12686
rect 56252 10780 56308 10836
rect 56364 11228 56420 11284
rect 55468 10332 55524 10388
rect 55020 7980 55076 8036
rect 55244 9996 55300 10052
rect 55356 9042 55412 9044
rect 55356 8990 55358 9042
rect 55358 8990 55410 9042
rect 55410 8990 55412 9042
rect 55356 8988 55412 8990
rect 51286 5514 51342 5516
rect 49532 5292 49588 5348
rect 50876 5404 50932 5460
rect 51286 5462 51288 5514
rect 51288 5462 51340 5514
rect 51340 5462 51342 5514
rect 51286 5460 51342 5462
rect 51390 5514 51446 5516
rect 51390 5462 51392 5514
rect 51392 5462 51444 5514
rect 51444 5462 51446 5514
rect 51390 5460 51446 5462
rect 51494 5514 51550 5516
rect 51494 5462 51496 5514
rect 51496 5462 51548 5514
rect 51548 5462 51550 5514
rect 51494 5460 51550 5462
rect 49756 5234 49812 5236
rect 49756 5182 49758 5234
rect 49758 5182 49810 5234
rect 49810 5182 49812 5234
rect 49756 5180 49812 5182
rect 51324 5292 51380 5348
rect 51100 5068 51156 5124
rect 48972 4844 49028 4900
rect 49644 4898 49700 4900
rect 49644 4846 49646 4898
rect 49646 4846 49698 4898
rect 49698 4846 49700 4898
rect 49644 4844 49700 4846
rect 49868 4508 49924 4564
rect 48860 4396 48916 4452
rect 49308 4396 49364 4452
rect 54012 5740 54068 5796
rect 53900 5404 53956 5460
rect 57484 12348 57540 12404
rect 57708 12290 57764 12292
rect 57708 12238 57710 12290
rect 57710 12238 57762 12290
rect 57762 12238 57764 12290
rect 57708 12236 57764 12238
rect 57260 11788 57316 11844
rect 57148 11228 57204 11284
rect 58439 14138 58495 14140
rect 58439 14086 58441 14138
rect 58441 14086 58493 14138
rect 58493 14086 58495 14138
rect 58439 14084 58495 14086
rect 58543 14138 58599 14140
rect 58543 14086 58545 14138
rect 58545 14086 58597 14138
rect 58597 14086 58599 14138
rect 58543 14084 58599 14086
rect 58647 14138 58703 14140
rect 58647 14086 58649 14138
rect 58649 14086 58701 14138
rect 58701 14086 58703 14138
rect 58647 14084 58703 14086
rect 58044 13356 58100 13412
rect 57932 12850 57988 12852
rect 57932 12798 57934 12850
rect 57934 12798 57986 12850
rect 57986 12798 57988 12850
rect 57932 12796 57988 12798
rect 57932 12178 57988 12180
rect 57932 12126 57934 12178
rect 57934 12126 57986 12178
rect 57986 12126 57988 12178
rect 57932 12124 57988 12126
rect 58439 12570 58495 12572
rect 58439 12518 58441 12570
rect 58441 12518 58493 12570
rect 58493 12518 58495 12570
rect 58439 12516 58495 12518
rect 58543 12570 58599 12572
rect 58543 12518 58545 12570
rect 58545 12518 58597 12570
rect 58597 12518 58599 12570
rect 58543 12516 58599 12518
rect 58647 12570 58703 12572
rect 58647 12518 58649 12570
rect 58649 12518 58701 12570
rect 58701 12518 58703 12570
rect 58647 12516 58703 12518
rect 58156 12348 58212 12404
rect 58156 12012 58212 12068
rect 57596 11788 57652 11844
rect 57820 11676 57876 11732
rect 57372 11170 57428 11172
rect 57372 11118 57374 11170
rect 57374 11118 57426 11170
rect 57426 11118 57428 11170
rect 57372 11116 57428 11118
rect 56924 10610 56980 10612
rect 56924 10558 56926 10610
rect 56926 10558 56978 10610
rect 56978 10558 56980 10610
rect 56924 10556 56980 10558
rect 56700 9996 56756 10052
rect 57372 9660 57428 9716
rect 58439 11002 58495 11004
rect 58439 10950 58441 11002
rect 58441 10950 58493 11002
rect 58493 10950 58495 11002
rect 58439 10948 58495 10950
rect 58543 11002 58599 11004
rect 58543 10950 58545 11002
rect 58545 10950 58597 11002
rect 58597 10950 58599 11002
rect 58543 10948 58599 10950
rect 58647 11002 58703 11004
rect 58647 10950 58649 11002
rect 58649 10950 58701 11002
rect 58701 10950 58703 11002
rect 58647 10948 58703 10950
rect 57932 10108 57988 10164
rect 56476 8428 56532 8484
rect 55580 8204 55636 8260
rect 55468 5794 55524 5796
rect 55468 5742 55470 5794
rect 55470 5742 55522 5794
rect 55522 5742 55524 5794
rect 55468 5740 55524 5742
rect 55356 5628 55412 5684
rect 57036 7532 57092 7588
rect 56140 6636 56196 6692
rect 55692 5964 55748 6020
rect 55692 5516 55748 5572
rect 54348 5292 54404 5348
rect 55356 5404 55412 5460
rect 52220 5068 52276 5124
rect 54572 5122 54628 5124
rect 54572 5070 54574 5122
rect 54574 5070 54626 5122
rect 54626 5070 54628 5122
rect 54572 5068 54628 5070
rect 55804 5292 55860 5348
rect 55692 5180 55748 5236
rect 51548 4450 51604 4452
rect 51548 4398 51550 4450
rect 51550 4398 51602 4450
rect 51602 4398 51604 4450
rect 51548 4396 51604 4398
rect 49532 4172 49588 4228
rect 51286 3946 51342 3948
rect 51286 3894 51288 3946
rect 51288 3894 51340 3946
rect 51340 3894 51342 3946
rect 51286 3892 51342 3894
rect 51390 3946 51446 3948
rect 51390 3894 51392 3946
rect 51392 3894 51444 3946
rect 51444 3894 51446 3946
rect 51390 3892 51446 3894
rect 51494 3946 51550 3948
rect 51494 3894 51496 3946
rect 51496 3894 51548 3946
rect 51548 3894 51550 3946
rect 51494 3892 51550 3894
rect 55804 5068 55860 5124
rect 56028 5180 56084 5236
rect 57148 7474 57204 7476
rect 57148 7422 57150 7474
rect 57150 7422 57202 7474
rect 57202 7422 57204 7474
rect 57148 7420 57204 7422
rect 57148 6860 57204 6916
rect 56924 5906 56980 5908
rect 56924 5854 56926 5906
rect 56926 5854 56978 5906
rect 56978 5854 56980 5906
rect 56924 5852 56980 5854
rect 56812 5180 56868 5236
rect 56588 5068 56644 5124
rect 55916 4226 55972 4228
rect 55916 4174 55918 4226
rect 55918 4174 55970 4226
rect 55970 4174 55972 4226
rect 55916 4172 55972 4174
rect 57596 7532 57652 7588
rect 57372 6690 57428 6692
rect 57372 6638 57374 6690
rect 57374 6638 57426 6690
rect 57426 6638 57428 6690
rect 57372 6636 57428 6638
rect 57260 5964 57316 6020
rect 56924 4396 56980 4452
rect 57036 5404 57092 5460
rect 1820 3276 1876 3332
rect 15518 3162 15574 3164
rect 15518 3110 15520 3162
rect 15520 3110 15572 3162
rect 15572 3110 15574 3162
rect 15518 3108 15574 3110
rect 15622 3162 15678 3164
rect 15622 3110 15624 3162
rect 15624 3110 15676 3162
rect 15676 3110 15678 3162
rect 15622 3108 15678 3110
rect 15726 3162 15782 3164
rect 15726 3110 15728 3162
rect 15728 3110 15780 3162
rect 15780 3110 15782 3162
rect 15726 3108 15782 3110
rect 29825 3162 29881 3164
rect 29825 3110 29827 3162
rect 29827 3110 29879 3162
rect 29879 3110 29881 3162
rect 29825 3108 29881 3110
rect 29929 3162 29985 3164
rect 29929 3110 29931 3162
rect 29931 3110 29983 3162
rect 29983 3110 29985 3162
rect 29929 3108 29985 3110
rect 30033 3162 30089 3164
rect 30033 3110 30035 3162
rect 30035 3110 30087 3162
rect 30087 3110 30089 3162
rect 30033 3108 30089 3110
rect 44132 3162 44188 3164
rect 44132 3110 44134 3162
rect 44134 3110 44186 3162
rect 44186 3110 44188 3162
rect 44132 3108 44188 3110
rect 44236 3162 44292 3164
rect 44236 3110 44238 3162
rect 44238 3110 44290 3162
rect 44290 3110 44292 3162
rect 44236 3108 44292 3110
rect 44340 3162 44396 3164
rect 44340 3110 44342 3162
rect 44342 3110 44394 3162
rect 44394 3110 44396 3162
rect 44340 3108 44396 3110
rect 57596 5740 57652 5796
rect 57484 5122 57540 5124
rect 57484 5070 57486 5122
rect 57486 5070 57538 5122
rect 57538 5070 57540 5122
rect 57484 5068 57540 5070
rect 58044 7474 58100 7476
rect 58044 7422 58046 7474
rect 58046 7422 58098 7474
rect 58098 7422 58100 7474
rect 58044 7420 58100 7422
rect 57820 5628 57876 5684
rect 57708 5404 57764 5460
rect 58044 5906 58100 5908
rect 58044 5854 58046 5906
rect 58046 5854 58098 5906
rect 58098 5854 58100 5906
rect 58044 5852 58100 5854
rect 57932 5068 57988 5124
rect 58439 9434 58495 9436
rect 58439 9382 58441 9434
rect 58441 9382 58493 9434
rect 58493 9382 58495 9434
rect 58439 9380 58495 9382
rect 58543 9434 58599 9436
rect 58543 9382 58545 9434
rect 58545 9382 58597 9434
rect 58597 9382 58599 9434
rect 58543 9380 58599 9382
rect 58647 9434 58703 9436
rect 58647 9382 58649 9434
rect 58649 9382 58701 9434
rect 58701 9382 58703 9434
rect 58647 9380 58703 9382
rect 58439 7866 58495 7868
rect 58439 7814 58441 7866
rect 58441 7814 58493 7866
rect 58493 7814 58495 7866
rect 58439 7812 58495 7814
rect 58543 7866 58599 7868
rect 58543 7814 58545 7866
rect 58545 7814 58597 7866
rect 58597 7814 58599 7866
rect 58543 7812 58599 7814
rect 58647 7866 58703 7868
rect 58647 7814 58649 7866
rect 58649 7814 58701 7866
rect 58701 7814 58703 7866
rect 58647 7812 58703 7814
rect 58439 6298 58495 6300
rect 58439 6246 58441 6298
rect 58441 6246 58493 6298
rect 58493 6246 58495 6298
rect 58439 6244 58495 6246
rect 58543 6298 58599 6300
rect 58543 6246 58545 6298
rect 58545 6246 58597 6298
rect 58597 6246 58599 6298
rect 58543 6244 58599 6246
rect 58647 6298 58703 6300
rect 58647 6246 58649 6298
rect 58649 6246 58701 6298
rect 58701 6246 58703 6298
rect 58647 6244 58703 6246
rect 58439 4730 58495 4732
rect 58439 4678 58441 4730
rect 58441 4678 58493 4730
rect 58493 4678 58495 4730
rect 58439 4676 58495 4678
rect 58543 4730 58599 4732
rect 58543 4678 58545 4730
rect 58545 4678 58597 4730
rect 58597 4678 58599 4730
rect 58543 4676 58599 4678
rect 58647 4730 58703 4732
rect 58647 4678 58649 4730
rect 58649 4678 58701 4730
rect 58701 4678 58703 4730
rect 58647 4676 58703 4678
rect 57932 4172 57988 4228
rect 58439 3162 58495 3164
rect 58439 3110 58441 3162
rect 58441 3110 58493 3162
rect 58493 3110 58495 3162
rect 58439 3108 58495 3110
rect 58543 3162 58599 3164
rect 58543 3110 58545 3162
rect 58545 3110 58597 3162
rect 58597 3110 58599 3162
rect 58543 3108 58599 3110
rect 58647 3162 58703 3164
rect 58647 3110 58649 3162
rect 58649 3110 58701 3162
rect 58701 3110 58703 3162
rect 58647 3108 58703 3110
rect 56252 2940 56308 2996
rect 1708 1372 1764 1428
<< metal3 >>
rect 0 28308 800 28336
rect 0 28252 5516 28308
rect 5572 28252 5582 28308
rect 0 28224 800 28252
rect 59200 27412 60000 27440
rect 57698 27356 57708 27412
rect 57764 27356 60000 27412
rect 59200 27328 60000 27356
rect 15508 26628 15518 26684
rect 15574 26628 15622 26684
rect 15678 26628 15726 26684
rect 15782 26628 15792 26684
rect 29815 26628 29825 26684
rect 29881 26628 29929 26684
rect 29985 26628 30033 26684
rect 30089 26628 30099 26684
rect 44122 26628 44132 26684
rect 44188 26628 44236 26684
rect 44292 26628 44340 26684
rect 44396 26628 44406 26684
rect 58429 26628 58439 26684
rect 58495 26628 58543 26684
rect 58599 26628 58647 26684
rect 58703 26628 58713 26684
rect 0 26516 800 26544
rect 0 26460 2156 26516
rect 2212 26460 2222 26516
rect 7970 26460 7980 26516
rect 8036 26460 13580 26516
rect 13636 26460 13646 26516
rect 21298 26460 21308 26516
rect 21364 26460 26684 26516
rect 26740 26460 26750 26516
rect 26852 26460 31332 26516
rect 50306 26460 50316 26516
rect 50372 26460 52220 26516
rect 52276 26460 52286 26516
rect 0 26432 800 26460
rect 1474 26348 1484 26404
rect 1540 26348 9324 26404
rect 9380 26348 9884 26404
rect 9940 26348 9950 26404
rect 15092 26348 16044 26404
rect 16100 26348 16110 26404
rect 16370 26348 16380 26404
rect 16436 26348 20748 26404
rect 20804 26348 21532 26404
rect 21588 26348 22092 26404
rect 22148 26348 22158 26404
rect 7298 26236 7308 26292
rect 7364 26236 10220 26292
rect 10276 26236 11340 26292
rect 11396 26236 11406 26292
rect 15092 26180 15148 26348
rect 26852 26292 26908 26460
rect 28914 26348 28924 26404
rect 28980 26348 29932 26404
rect 29988 26348 29998 26404
rect 31276 26292 31332 26460
rect 36082 26348 36092 26404
rect 36148 26348 39116 26404
rect 39172 26348 40124 26404
rect 40180 26348 40190 26404
rect 16258 26236 16268 26292
rect 16324 26236 17500 26292
rect 17556 26236 17566 26292
rect 22642 26236 22652 26292
rect 22708 26236 26908 26292
rect 26964 26236 26974 26292
rect 27346 26236 27356 26292
rect 27412 26236 28700 26292
rect 28756 26236 28766 26292
rect 31266 26236 31276 26292
rect 31332 26236 31342 26292
rect 35522 26236 35532 26292
rect 35588 26236 36204 26292
rect 36260 26236 36270 26292
rect 49522 26236 49532 26292
rect 49588 26236 49598 26292
rect 49970 26236 49980 26292
rect 50036 26236 50428 26292
rect 50484 26236 50494 26292
rect 49532 26180 49588 26236
rect 3332 26124 5964 26180
rect 6020 26124 6030 26180
rect 8866 26124 8876 26180
rect 8932 26124 15148 26180
rect 19618 26124 19628 26180
rect 19684 26124 21084 26180
rect 21140 26124 21150 26180
rect 24658 26124 24668 26180
rect 24724 26124 25452 26180
rect 25508 26124 26908 26180
rect 34178 26124 34188 26180
rect 34244 26124 35420 26180
rect 35476 26124 35486 26180
rect 35970 26124 35980 26180
rect 36036 26124 39900 26180
rect 39956 26124 39966 26180
rect 40226 26124 40236 26180
rect 40292 26124 46844 26180
rect 46900 26124 48076 26180
rect 48132 26124 48636 26180
rect 48692 26124 48702 26180
rect 49532 26124 51772 26180
rect 51828 26124 51838 26180
rect 3332 26068 3388 26124
rect 1250 26012 1260 26068
rect 1316 26012 3388 26068
rect 7634 26012 7644 26068
rect 7700 26012 11116 26068
rect 11172 26012 11182 26068
rect 15026 26012 15036 26068
rect 15092 26012 19180 26068
rect 19236 26012 19964 26068
rect 20020 26012 20030 26068
rect 22082 26012 22092 26068
rect 22148 26012 23660 26068
rect 23716 26012 23726 26068
rect 23986 26012 23996 26068
rect 24052 26012 25228 26068
rect 25284 26012 25294 26068
rect 26852 25956 26908 26124
rect 35420 26068 35476 26124
rect 35420 26012 37436 26068
rect 37492 26012 37502 26068
rect 49186 26012 49196 26068
rect 49252 26012 50204 26068
rect 50260 26012 50270 26068
rect 50418 26012 50428 26068
rect 50484 26012 51212 26068
rect 51268 26012 51278 26068
rect 26852 25900 27020 25956
rect 27076 25900 31948 25956
rect 32004 25900 32014 25956
rect 8355 25844 8365 25900
rect 8421 25844 8469 25900
rect 8525 25844 8573 25900
rect 8629 25844 8639 25900
rect 22662 25844 22672 25900
rect 22728 25844 22776 25900
rect 22832 25844 22880 25900
rect 22936 25844 22946 25900
rect 36969 25844 36979 25900
rect 37035 25844 37083 25900
rect 37139 25844 37187 25900
rect 37243 25844 37253 25900
rect 51276 25844 51286 25900
rect 51342 25844 51390 25900
rect 51446 25844 51494 25900
rect 51550 25844 51560 25900
rect 8754 25788 8764 25844
rect 8820 25788 9772 25844
rect 9828 25788 20076 25844
rect 20132 25788 20142 25844
rect 23090 25788 23100 25844
rect 23156 25788 26012 25844
rect 26068 25788 26078 25844
rect 26226 25788 26236 25844
rect 26292 25788 27356 25844
rect 27412 25788 27422 25844
rect 8764 25732 8820 25788
rect 4050 25676 4060 25732
rect 4116 25676 5852 25732
rect 5908 25676 7196 25732
rect 7252 25676 8820 25732
rect 9874 25676 9884 25732
rect 9940 25676 47628 25732
rect 47684 25676 47694 25732
rect 6850 25564 6860 25620
rect 6916 25564 7532 25620
rect 7588 25564 9436 25620
rect 9492 25564 9502 25620
rect 12002 25564 12012 25620
rect 12068 25564 13244 25620
rect 13300 25564 14364 25620
rect 14420 25564 14430 25620
rect 26450 25564 26460 25620
rect 26516 25564 29372 25620
rect 29428 25564 29820 25620
rect 29876 25564 31612 25620
rect 31668 25564 32396 25620
rect 32452 25564 35532 25620
rect 35588 25564 35598 25620
rect 36204 25564 38668 25620
rect 47506 25564 47516 25620
rect 47572 25564 56588 25620
rect 56644 25564 56654 25620
rect 36204 25508 36260 25564
rect 38612 25508 38668 25564
rect 3332 25452 8092 25508
rect 8148 25452 8158 25508
rect 11890 25452 11900 25508
rect 11956 25452 12460 25508
rect 12516 25452 13468 25508
rect 13524 25452 13534 25508
rect 14466 25452 14476 25508
rect 14532 25452 15148 25508
rect 15204 25452 15214 25508
rect 17602 25452 17612 25508
rect 17668 25452 19068 25508
rect 19124 25452 19134 25508
rect 32050 25452 32060 25508
rect 32116 25452 32732 25508
rect 32788 25452 32798 25508
rect 36194 25452 36204 25508
rect 36260 25452 36270 25508
rect 36418 25452 36428 25508
rect 36484 25452 37548 25508
rect 37604 25452 37614 25508
rect 38612 25452 38780 25508
rect 38836 25452 38846 25508
rect 52994 25452 53004 25508
rect 53060 25452 53676 25508
rect 53732 25452 55468 25508
rect 55524 25452 55534 25508
rect 3332 25396 3388 25452
rect 3042 25340 3052 25396
rect 3108 25340 3388 25396
rect 6962 25340 6972 25396
rect 7028 25340 9100 25396
rect 9156 25340 9166 25396
rect 9762 25340 9772 25396
rect 9828 25340 16268 25396
rect 16324 25340 16334 25396
rect 16706 25340 16716 25396
rect 16772 25340 18732 25396
rect 18788 25340 18798 25396
rect 19730 25340 19740 25396
rect 19796 25340 20972 25396
rect 21028 25340 21308 25396
rect 21364 25340 21374 25396
rect 28466 25340 28476 25396
rect 28532 25340 32844 25396
rect 32900 25340 32910 25396
rect 35410 25340 35420 25396
rect 35476 25340 41356 25396
rect 41412 25340 41422 25396
rect 42690 25340 42700 25396
rect 42756 25340 44492 25396
rect 44548 25340 45276 25396
rect 45332 25340 45342 25396
rect 47842 25340 47852 25396
rect 47908 25340 49196 25396
rect 49252 25340 49262 25396
rect 4834 25228 4844 25284
rect 4900 25228 7644 25284
rect 7700 25228 7710 25284
rect 11442 25228 11452 25284
rect 11508 25228 12348 25284
rect 12404 25228 12414 25284
rect 16482 25228 16492 25284
rect 16548 25228 18060 25284
rect 18116 25228 18126 25284
rect 34962 25228 34972 25284
rect 35028 25228 35812 25284
rect 36306 25228 36316 25284
rect 36372 25228 44716 25284
rect 44772 25228 45164 25284
rect 45220 25228 45230 25284
rect 48178 25228 48188 25284
rect 48244 25228 48972 25284
rect 49028 25228 49038 25284
rect 35756 25172 35812 25228
rect 31154 25116 31164 25172
rect 31220 25116 31836 25172
rect 31892 25116 33740 25172
rect 33796 25116 33806 25172
rect 35746 25116 35756 25172
rect 35812 25116 37436 25172
rect 37492 25116 37996 25172
rect 38052 25116 38062 25172
rect 15508 25060 15518 25116
rect 15574 25060 15622 25116
rect 15678 25060 15726 25116
rect 15782 25060 15792 25116
rect 29815 25060 29825 25116
rect 29881 25060 29929 25116
rect 29985 25060 30033 25116
rect 30089 25060 30099 25116
rect 44122 25060 44132 25116
rect 44188 25060 44236 25116
rect 44292 25060 44340 25116
rect 44396 25060 44406 25116
rect 58429 25060 58439 25116
rect 58495 25060 58543 25116
rect 58599 25060 58647 25116
rect 58703 25060 58713 25116
rect 7186 25004 7196 25060
rect 7252 25004 8988 25060
rect 9044 25004 9054 25060
rect 31714 25004 31724 25060
rect 31780 25004 40236 25060
rect 40292 25004 40302 25060
rect 29586 24892 29596 24948
rect 29652 24892 30604 24948
rect 30660 24892 31388 24948
rect 31444 24892 31454 24948
rect 34962 24892 34972 24948
rect 35028 24892 36988 24948
rect 37044 24892 37054 24948
rect 5618 24780 5628 24836
rect 5684 24780 15148 24836
rect 23426 24780 23436 24836
rect 23492 24780 24668 24836
rect 24724 24780 26908 24836
rect 31042 24780 31052 24836
rect 31108 24780 32172 24836
rect 32228 24780 32238 24836
rect 32386 24780 32396 24836
rect 32452 24780 33404 24836
rect 33460 24780 34188 24836
rect 34244 24780 34748 24836
rect 34804 24780 34814 24836
rect 36418 24780 36428 24836
rect 36484 24780 37212 24836
rect 37268 24780 37278 24836
rect 0 24724 800 24752
rect 0 24668 1708 24724
rect 1764 24668 4732 24724
rect 4788 24668 4798 24724
rect 6626 24668 6636 24724
rect 6692 24668 10892 24724
rect 10948 24668 12236 24724
rect 12292 24668 12302 24724
rect 12562 24668 12572 24724
rect 12628 24668 13356 24724
rect 13412 24668 13422 24724
rect 15092 24668 15148 24780
rect 26852 24724 26908 24780
rect 15204 24668 15214 24724
rect 16034 24668 16044 24724
rect 16100 24668 18396 24724
rect 18452 24668 18462 24724
rect 20626 24668 20636 24724
rect 20692 24668 22540 24724
rect 22596 24668 22606 24724
rect 26852 24668 28364 24724
rect 28420 24668 29596 24724
rect 29652 24668 30492 24724
rect 30548 24668 30558 24724
rect 31378 24668 31388 24724
rect 31444 24668 33180 24724
rect 33236 24668 33246 24724
rect 33506 24668 33516 24724
rect 33572 24668 39564 24724
rect 39620 24668 41692 24724
rect 41748 24668 41758 24724
rect 42690 24668 42700 24724
rect 42756 24668 45948 24724
rect 46004 24668 46508 24724
rect 46564 24668 46574 24724
rect 0 24640 800 24668
rect 9874 24556 9884 24612
rect 9940 24556 13468 24612
rect 13524 24556 13534 24612
rect 21186 24556 21196 24612
rect 21252 24556 21644 24612
rect 21700 24556 22204 24612
rect 22260 24556 22270 24612
rect 42242 24556 42252 24612
rect 42308 24556 42924 24612
rect 42980 24556 42990 24612
rect 43250 24556 43260 24612
rect 43316 24556 48188 24612
rect 48244 24556 50540 24612
rect 50596 24556 50606 24612
rect 6626 24444 6636 24500
rect 6692 24444 7756 24500
rect 7812 24444 7822 24500
rect 15698 24444 15708 24500
rect 15764 24444 17500 24500
rect 17556 24444 17566 24500
rect 22428 24444 22652 24500
rect 22708 24444 24444 24500
rect 24500 24444 25340 24500
rect 25396 24444 25406 24500
rect 22428 24388 22484 24444
rect 16818 24332 16828 24388
rect 16884 24332 20412 24388
rect 20468 24332 21980 24388
rect 22036 24332 22046 24388
rect 22418 24332 22428 24388
rect 22484 24332 22494 24388
rect 8355 24276 8365 24332
rect 8421 24276 8469 24332
rect 8525 24276 8573 24332
rect 8629 24276 8639 24332
rect 22662 24276 22672 24332
rect 22728 24276 22776 24332
rect 22832 24276 22880 24332
rect 22936 24276 22946 24332
rect 36969 24276 36979 24332
rect 37035 24276 37083 24332
rect 37139 24276 37187 24332
rect 37243 24276 37253 24332
rect 51276 24276 51286 24332
rect 51342 24276 51390 24332
rect 51446 24276 51494 24332
rect 51550 24276 51560 24332
rect 13458 24220 13468 24276
rect 13524 24220 18508 24276
rect 18564 24220 18574 24276
rect 21858 24220 21868 24276
rect 21924 24220 22316 24276
rect 22372 24220 22382 24276
rect 8194 24108 8204 24164
rect 8260 24108 8876 24164
rect 8932 24108 10220 24164
rect 10276 24108 11004 24164
rect 11060 24108 14028 24164
rect 14084 24108 14094 24164
rect 15092 24108 16156 24164
rect 16212 24108 16222 24164
rect 22194 24108 22204 24164
rect 22260 24108 22764 24164
rect 22820 24108 22830 24164
rect 33170 24108 33180 24164
rect 33236 24108 34524 24164
rect 34580 24108 34590 24164
rect 15092 24052 15148 24108
rect 3266 23996 3276 24052
rect 3332 23996 6412 24052
rect 6468 23996 6478 24052
rect 7186 23996 7196 24052
rect 7252 23996 12236 24052
rect 12292 23996 12302 24052
rect 12898 23996 12908 24052
rect 12964 23996 15148 24052
rect 20066 23996 20076 24052
rect 20132 23996 26236 24052
rect 26292 23996 26908 24052
rect 34738 23996 34748 24052
rect 34804 23996 35420 24052
rect 35476 23996 35486 24052
rect 8978 23884 8988 23940
rect 9044 23884 10332 23940
rect 10388 23884 11900 23940
rect 11956 23884 11966 23940
rect 13346 23884 13356 23940
rect 13412 23884 14028 23940
rect 14084 23884 14476 23940
rect 14532 23884 14542 23940
rect 17266 23884 17276 23940
rect 17332 23884 17948 23940
rect 18004 23884 19964 23940
rect 20020 23884 20030 23940
rect 13356 23828 13412 23884
rect 26852 23828 26908 23996
rect 27794 23884 27804 23940
rect 27860 23884 28588 23940
rect 28644 23884 28654 23940
rect 35858 23884 35868 23940
rect 35924 23884 39228 23940
rect 39284 23884 39294 23940
rect 46834 23884 46844 23940
rect 46900 23884 48636 23940
rect 48692 23884 50428 23940
rect 54898 23884 54908 23940
rect 54964 23884 55580 23940
rect 55636 23884 57708 23940
rect 57764 23884 57774 23940
rect 50372 23828 50428 23884
rect 59200 23828 60000 23856
rect 4610 23772 4620 23828
rect 4676 23772 5180 23828
rect 5236 23772 7196 23828
rect 7252 23772 7262 23828
rect 8306 23772 8316 23828
rect 8372 23772 13412 23828
rect 16034 23772 16044 23828
rect 16100 23772 20636 23828
rect 20692 23772 21980 23828
rect 22036 23772 22046 23828
rect 22194 23772 22204 23828
rect 22260 23772 22540 23828
rect 22596 23772 24780 23828
rect 24836 23772 24846 23828
rect 26852 23772 29260 23828
rect 29316 23772 29326 23828
rect 39330 23772 39340 23828
rect 39396 23772 41020 23828
rect 41076 23772 42140 23828
rect 42196 23772 42206 23828
rect 44482 23772 44492 23828
rect 44548 23772 47180 23828
rect 47236 23772 48748 23828
rect 48804 23772 48814 23828
rect 50372 23772 51324 23828
rect 51380 23772 51884 23828
rect 51940 23772 51950 23828
rect 52882 23772 52892 23828
rect 52948 23772 52958 23828
rect 57596 23772 60000 23828
rect 52892 23716 52948 23772
rect 57596 23716 57652 23772
rect 59200 23744 60000 23772
rect 6626 23660 6636 23716
rect 6692 23660 10780 23716
rect 10836 23660 10846 23716
rect 15250 23660 15260 23716
rect 15316 23660 22428 23716
rect 22484 23660 22494 23716
rect 26674 23660 26684 23716
rect 26740 23660 28700 23716
rect 28756 23660 28766 23716
rect 33394 23660 33404 23716
rect 33460 23660 35308 23716
rect 35364 23660 36428 23716
rect 36484 23660 36494 23716
rect 52210 23660 52220 23716
rect 52276 23660 53564 23716
rect 53620 23660 53630 23716
rect 57586 23660 57596 23716
rect 57652 23660 57662 23716
rect 12226 23548 12236 23604
rect 12292 23548 13580 23604
rect 13636 23548 13646 23604
rect 18386 23548 18396 23604
rect 18452 23548 22540 23604
rect 22596 23548 22606 23604
rect 25778 23548 25788 23604
rect 25844 23548 29148 23604
rect 29204 23548 29214 23604
rect 38098 23548 38108 23604
rect 38164 23548 39116 23604
rect 39172 23548 39182 23604
rect 40562 23548 40572 23604
rect 40628 23548 43260 23604
rect 43316 23548 43326 23604
rect 54562 23548 54572 23604
rect 54628 23548 57932 23604
rect 57988 23548 57998 23604
rect 15508 23492 15518 23548
rect 15574 23492 15622 23548
rect 15678 23492 15726 23548
rect 15782 23492 15792 23548
rect 29815 23492 29825 23548
rect 29881 23492 29929 23548
rect 29985 23492 30033 23548
rect 30089 23492 30099 23548
rect 44122 23492 44132 23548
rect 44188 23492 44236 23548
rect 44292 23492 44340 23548
rect 44396 23492 44406 23548
rect 58429 23492 58439 23548
rect 58495 23492 58543 23548
rect 58599 23492 58647 23548
rect 58703 23492 58713 23548
rect 2146 23436 2156 23492
rect 2212 23436 7532 23492
rect 7588 23436 7598 23492
rect 20188 23436 21868 23492
rect 21924 23436 23324 23492
rect 23380 23436 23390 23492
rect 24434 23436 24444 23492
rect 24500 23436 26348 23492
rect 26404 23436 27132 23492
rect 27188 23436 27198 23492
rect 30370 23436 30380 23492
rect 30436 23436 31948 23492
rect 32004 23436 32014 23492
rect 20188 23380 20244 23436
rect 11666 23324 11676 23380
rect 11732 23324 16716 23380
rect 16772 23324 16782 23380
rect 16930 23324 16940 23380
rect 16996 23324 20188 23380
rect 20244 23324 20254 23380
rect 21410 23324 21420 23380
rect 21476 23324 22316 23380
rect 22372 23324 22382 23380
rect 24546 23324 24556 23380
rect 24612 23324 25676 23380
rect 25732 23324 27020 23380
rect 27076 23324 31052 23380
rect 31108 23324 31118 23380
rect 38612 23324 39676 23380
rect 39732 23324 39742 23380
rect 52658 23324 52668 23380
rect 52724 23324 55804 23380
rect 55860 23324 57036 23380
rect 57092 23324 57102 23380
rect 2930 23212 2940 23268
rect 2996 23212 3724 23268
rect 3780 23212 3790 23268
rect 4722 23212 4732 23268
rect 4788 23212 13132 23268
rect 13188 23212 13198 23268
rect 18050 23212 18060 23268
rect 18116 23212 21532 23268
rect 21588 23212 21598 23268
rect 26852 23212 35812 23268
rect 26852 23156 26908 23212
rect 35756 23156 35812 23212
rect 38612 23156 38668 23324
rect 49522 23212 49532 23268
rect 49588 23212 49756 23268
rect 49812 23212 49822 23268
rect 52098 23212 52108 23268
rect 52164 23212 52444 23268
rect 52500 23212 53228 23268
rect 53284 23212 53294 23268
rect 55458 23212 55468 23268
rect 55524 23212 56924 23268
rect 56980 23212 56990 23268
rect 2258 23100 2268 23156
rect 2324 23100 3836 23156
rect 3892 23100 4620 23156
rect 4676 23100 4686 23156
rect 5394 23100 5404 23156
rect 5460 23100 9100 23156
rect 9156 23100 9772 23156
rect 9828 23100 9838 23156
rect 11890 23100 11900 23156
rect 11956 23100 12684 23156
rect 12740 23100 12750 23156
rect 23874 23100 23884 23156
rect 23940 23100 26908 23156
rect 29698 23100 29708 23156
rect 29764 23100 33740 23156
rect 33796 23100 34412 23156
rect 34468 23100 35308 23156
rect 35364 23100 35374 23156
rect 35746 23100 35756 23156
rect 35812 23100 35822 23156
rect 36866 23100 36876 23156
rect 36932 23100 38668 23156
rect 40338 23100 40348 23156
rect 40404 23100 41244 23156
rect 41300 23100 42028 23156
rect 42084 23100 42094 23156
rect 42242 23100 42252 23156
rect 42308 23100 42924 23156
rect 42980 23100 42990 23156
rect 47058 23100 47068 23156
rect 47124 23100 48412 23156
rect 48468 23100 48478 23156
rect 5058 22988 5068 23044
rect 5124 22988 6300 23044
rect 6356 22988 6366 23044
rect 16034 22988 16044 23044
rect 16100 22988 17836 23044
rect 17892 22988 17902 23044
rect 18274 22988 18284 23044
rect 18340 22988 25676 23044
rect 25732 22988 25742 23044
rect 26450 22988 26460 23044
rect 26516 22988 26526 23044
rect 0 22932 800 22960
rect 17836 22932 17892 22988
rect 26460 22932 26516 22988
rect 26852 22932 26908 23044
rect 26964 22988 26974 23044
rect 30482 22988 30492 23044
rect 30548 22988 31388 23044
rect 31444 22988 33628 23044
rect 33684 22988 33694 23044
rect 36306 22988 36316 23044
rect 36372 22988 37660 23044
rect 37716 22988 38108 23044
rect 38164 22988 38174 23044
rect 39890 22988 39900 23044
rect 39956 22988 43596 23044
rect 43652 22988 43662 23044
rect 0 22876 2604 22932
rect 2660 22876 4060 22932
rect 4116 22876 4126 22932
rect 4946 22876 4956 22932
rect 5012 22876 8876 22932
rect 8932 22876 8942 22932
rect 17836 22876 18620 22932
rect 18676 22876 18686 22932
rect 26460 22876 26908 22932
rect 28914 22876 28924 22932
rect 28980 22876 30380 22932
rect 30436 22876 30446 22932
rect 35074 22876 35084 22932
rect 35140 22876 35980 22932
rect 36036 22876 36046 22932
rect 37202 22876 37212 22932
rect 37268 22876 38612 22932
rect 0 22848 800 22876
rect 38556 22820 38612 22876
rect 50428 22876 52332 22932
rect 52388 22876 53004 22932
rect 53060 22876 53070 22932
rect 1810 22764 1820 22820
rect 1876 22764 2716 22820
rect 2772 22764 2782 22820
rect 5618 22764 5628 22820
rect 5684 22764 7308 22820
rect 7364 22764 7374 22820
rect 38546 22764 38556 22820
rect 38612 22764 41020 22820
rect 41076 22764 41086 22820
rect 8355 22708 8365 22764
rect 8421 22708 8469 22764
rect 8525 22708 8573 22764
rect 8629 22708 8639 22764
rect 22662 22708 22672 22764
rect 22728 22708 22776 22764
rect 22832 22708 22880 22764
rect 22936 22708 22946 22764
rect 36969 22708 36979 22764
rect 37035 22708 37083 22764
rect 37139 22708 37187 22764
rect 37243 22708 37253 22764
rect 50428 22708 50484 22876
rect 51276 22708 51286 22764
rect 51342 22708 51390 22764
rect 51446 22708 51494 22764
rect 51550 22708 51560 22764
rect 19618 22652 19628 22708
rect 19684 22652 20860 22708
rect 20916 22652 20926 22708
rect 24444 22652 25228 22708
rect 25284 22652 25294 22708
rect 26786 22652 26796 22708
rect 26852 22652 28028 22708
rect 28084 22652 28588 22708
rect 28644 22652 28654 22708
rect 38612 22652 50428 22708
rect 50484 22652 50494 22708
rect 24444 22596 24500 22652
rect 14130 22540 14140 22596
rect 14196 22540 15036 22596
rect 15092 22540 15102 22596
rect 16034 22540 16044 22596
rect 16100 22540 16940 22596
rect 16996 22540 17836 22596
rect 17892 22540 17902 22596
rect 21858 22540 21868 22596
rect 21924 22540 22988 22596
rect 23044 22540 24500 22596
rect 24658 22540 24668 22596
rect 24724 22540 36204 22596
rect 36260 22540 36270 22596
rect 38612 22484 38668 22652
rect 46946 22540 46956 22596
rect 47012 22540 52780 22596
rect 52836 22540 52846 22596
rect 8082 22428 8092 22484
rect 8148 22428 38668 22484
rect 39666 22428 39676 22484
rect 39732 22428 41468 22484
rect 41524 22428 41534 22484
rect 44258 22428 44268 22484
rect 44324 22428 46508 22484
rect 46564 22428 46574 22484
rect 48738 22428 48748 22484
rect 48804 22428 53004 22484
rect 53060 22428 53070 22484
rect 8866 22316 8876 22372
rect 8932 22316 13692 22372
rect 13748 22316 13758 22372
rect 15092 22316 16044 22372
rect 16100 22316 16110 22372
rect 16258 22316 16268 22372
rect 16324 22316 16362 22372
rect 22194 22316 22204 22372
rect 22260 22316 23548 22372
rect 23604 22316 23614 22372
rect 37538 22316 37548 22372
rect 37604 22316 38220 22372
rect 38276 22316 38286 22372
rect 38994 22316 39004 22372
rect 39060 22316 40012 22372
rect 40068 22316 40078 22372
rect 44818 22316 44828 22372
rect 44884 22316 47068 22372
rect 47124 22316 47134 22372
rect 47282 22316 47292 22372
rect 47348 22316 49532 22372
rect 49588 22316 49598 22372
rect 53330 22316 53340 22372
rect 53396 22316 53788 22372
rect 53844 22316 55132 22372
rect 55188 22316 56364 22372
rect 56420 22316 56430 22372
rect 15092 22260 15148 22316
rect 6290 22204 6300 22260
rect 6356 22204 8204 22260
rect 8260 22204 8270 22260
rect 13458 22204 13468 22260
rect 13524 22204 15148 22260
rect 22530 22204 22540 22260
rect 22596 22204 24332 22260
rect 24388 22204 24398 22260
rect 26786 22204 26796 22260
rect 26852 22204 36988 22260
rect 37044 22204 37054 22260
rect 45266 22204 45276 22260
rect 45332 22204 47964 22260
rect 48020 22204 49756 22260
rect 49812 22204 49822 22260
rect 53442 22204 53452 22260
rect 53508 22204 53676 22260
rect 53732 22204 54348 22260
rect 54404 22204 54414 22260
rect 13682 22092 13692 22148
rect 13748 22092 16268 22148
rect 16324 22092 16334 22148
rect 16594 22092 16604 22148
rect 16660 22092 18172 22148
rect 18228 22092 18238 22148
rect 20850 22092 20860 22148
rect 20916 22092 22764 22148
rect 22820 22092 22830 22148
rect 38546 22092 38556 22148
rect 38612 22092 41356 22148
rect 41412 22092 42364 22148
rect 42420 22092 42924 22148
rect 42980 22092 44044 22148
rect 44100 22092 44548 22148
rect 47730 22092 47740 22148
rect 47796 22092 52892 22148
rect 52948 22092 52958 22148
rect 44492 22036 44548 22092
rect 18386 21980 18396 22036
rect 18452 21980 22428 22036
rect 22484 21980 25676 22036
rect 25732 21980 25742 22036
rect 44492 21980 48972 22036
rect 49028 21980 49038 22036
rect 15508 21924 15518 21980
rect 15574 21924 15622 21980
rect 15678 21924 15726 21980
rect 15782 21924 15792 21980
rect 29815 21924 29825 21980
rect 29881 21924 29929 21980
rect 29985 21924 30033 21980
rect 30089 21924 30099 21980
rect 44122 21924 44132 21980
rect 44188 21924 44236 21980
rect 44292 21924 44340 21980
rect 44396 21924 44406 21980
rect 58429 21924 58439 21980
rect 58495 21924 58543 21980
rect 58599 21924 58647 21980
rect 58703 21924 58713 21980
rect 4946 21868 4956 21924
rect 5012 21868 11452 21924
rect 11508 21868 11676 21924
rect 11732 21868 11742 21924
rect 13010 21868 13020 21924
rect 13076 21868 13804 21924
rect 13860 21868 13870 21924
rect 46498 21868 46508 21924
rect 46564 21868 49532 21924
rect 49588 21868 49598 21924
rect 1698 21756 1708 21812
rect 1764 21756 2604 21812
rect 2660 21756 3388 21812
rect 3444 21756 3454 21812
rect 8866 21756 8876 21812
rect 8932 21756 14476 21812
rect 14532 21756 14542 21812
rect 16258 21756 16268 21812
rect 16324 21756 16604 21812
rect 16660 21756 16670 21812
rect 20738 21756 20748 21812
rect 20804 21756 21532 21812
rect 21588 21756 21598 21812
rect 26562 21756 26572 21812
rect 26628 21756 30380 21812
rect 30436 21756 34412 21812
rect 34468 21756 35308 21812
rect 35364 21756 35374 21812
rect 47618 21756 47628 21812
rect 47684 21756 49644 21812
rect 49700 21756 49710 21812
rect 51202 21756 51212 21812
rect 51268 21756 52052 21812
rect 54114 21756 54124 21812
rect 54180 21756 55356 21812
rect 55412 21756 55422 21812
rect 7410 21644 7420 21700
rect 7476 21644 10668 21700
rect 10724 21644 10734 21700
rect 13794 21644 13804 21700
rect 13860 21644 15148 21700
rect 21410 21644 21420 21700
rect 21476 21644 26124 21700
rect 26180 21644 26190 21700
rect 35410 21644 35420 21700
rect 35476 21644 36428 21700
rect 36484 21644 36494 21700
rect 45938 21644 45948 21700
rect 46004 21644 49308 21700
rect 49364 21644 49374 21700
rect 15092 21588 15148 21644
rect 51996 21588 52052 21756
rect 53554 21644 53564 21700
rect 53620 21644 55468 21700
rect 55524 21644 55534 21700
rect 3490 21532 3500 21588
rect 3556 21532 4508 21588
rect 4564 21532 4574 21588
rect 5170 21532 5180 21588
rect 5236 21532 6076 21588
rect 6132 21532 6142 21588
rect 8978 21532 8988 21588
rect 9044 21532 11564 21588
rect 11620 21532 11630 21588
rect 13906 21532 13916 21588
rect 13972 21532 13982 21588
rect 15092 21532 20412 21588
rect 20468 21532 22204 21588
rect 22260 21532 22270 21588
rect 23874 21532 23884 21588
rect 23940 21532 27020 21588
rect 27076 21532 27086 21588
rect 27682 21532 27692 21588
rect 27748 21532 31052 21588
rect 31108 21532 31118 21588
rect 37314 21532 37324 21588
rect 37380 21532 38332 21588
rect 38388 21532 38398 21588
rect 43586 21532 43596 21588
rect 43652 21532 48748 21588
rect 48804 21532 48814 21588
rect 51986 21532 51996 21588
rect 52052 21532 53900 21588
rect 53956 21532 54796 21588
rect 54852 21532 55244 21588
rect 55300 21532 55310 21588
rect 55794 21532 55804 21588
rect 55860 21532 57932 21588
rect 57988 21532 57998 21588
rect 5954 21420 5964 21476
rect 6020 21420 6300 21476
rect 6356 21420 6366 21476
rect 10546 21420 10556 21476
rect 10612 21420 10780 21476
rect 10836 21420 11900 21476
rect 11956 21420 11966 21476
rect 13916 21364 13972 21532
rect 55244 21476 55300 21532
rect 15922 21420 15932 21476
rect 15988 21420 17612 21476
rect 17668 21420 17678 21476
rect 20626 21420 20636 21476
rect 20692 21420 25676 21476
rect 25732 21420 25742 21476
rect 28466 21420 28476 21476
rect 28532 21420 28542 21476
rect 44034 21420 44044 21476
rect 44100 21420 46620 21476
rect 46676 21420 46686 21476
rect 47394 21420 47404 21476
rect 47460 21420 48188 21476
rect 48244 21420 48636 21476
rect 48692 21420 48702 21476
rect 55244 21420 56028 21476
rect 56084 21420 56700 21476
rect 56756 21420 56766 21476
rect 13916 21308 16044 21364
rect 16100 21308 16110 21364
rect 16258 21308 16268 21364
rect 16324 21308 16940 21364
rect 16996 21308 17006 21364
rect 28476 21252 28532 21420
rect 40226 21308 40236 21364
rect 40292 21308 42028 21364
rect 42084 21308 42094 21364
rect 23986 21196 23996 21252
rect 24052 21196 24556 21252
rect 24612 21196 30268 21252
rect 30324 21196 32396 21252
rect 32452 21196 34860 21252
rect 34916 21196 34926 21252
rect 0 21140 800 21168
rect 8355 21140 8365 21196
rect 8421 21140 8469 21196
rect 8525 21140 8573 21196
rect 8629 21140 8639 21196
rect 22662 21140 22672 21196
rect 22728 21140 22776 21196
rect 22832 21140 22880 21196
rect 22936 21140 22946 21196
rect 36969 21140 36979 21196
rect 37035 21140 37083 21196
rect 37139 21140 37187 21196
rect 37243 21140 37253 21196
rect 51276 21140 51286 21196
rect 51342 21140 51390 21196
rect 51446 21140 51494 21196
rect 51550 21140 51560 21196
rect 0 21084 1708 21140
rect 1764 21084 1820 21140
rect 1876 21084 1886 21140
rect 0 21056 800 21084
rect 6290 20972 6300 21028
rect 6356 20972 10892 21028
rect 10948 20972 10958 21028
rect 36418 20972 36428 21028
rect 36484 20972 36988 21028
rect 37044 20972 37054 21028
rect 42130 20972 42140 21028
rect 42196 20972 43708 21028
rect 43764 20972 47180 21028
rect 47236 20972 47246 21028
rect 50652 20972 52108 21028
rect 52164 20972 52174 21028
rect 50652 20916 50708 20972
rect 4498 20860 4508 20916
rect 4564 20860 5852 20916
rect 5908 20860 5918 20916
rect 6402 20860 6412 20916
rect 6468 20860 50652 20916
rect 50708 20860 50718 20916
rect 51874 20860 51884 20916
rect 51940 20860 54796 20916
rect 54852 20860 54862 20916
rect 4610 20748 4620 20804
rect 4676 20748 6748 20804
rect 6804 20748 6814 20804
rect 15250 20748 15260 20804
rect 15316 20748 16604 20804
rect 16660 20748 17052 20804
rect 17108 20748 17118 20804
rect 20738 20748 20748 20804
rect 20804 20748 22540 20804
rect 22596 20748 23324 20804
rect 23380 20748 23390 20804
rect 25330 20748 25340 20804
rect 25396 20748 28308 20804
rect 31602 20748 31612 20804
rect 31668 20748 31836 20804
rect 31892 20748 32172 20804
rect 32228 20748 32238 20804
rect 34514 20748 34524 20804
rect 34580 20748 38780 20804
rect 38836 20748 38846 20804
rect 42018 20748 42028 20804
rect 42084 20748 44492 20804
rect 44548 20748 46060 20804
rect 46116 20748 46126 20804
rect 46722 20748 46732 20804
rect 46788 20748 50764 20804
rect 50820 20748 50830 20804
rect 53442 20748 53452 20804
rect 53508 20748 55020 20804
rect 55076 20748 55086 20804
rect 28252 20692 28308 20748
rect 3266 20636 3276 20692
rect 3332 20636 4732 20692
rect 4788 20636 6860 20692
rect 6916 20636 6926 20692
rect 16034 20636 16044 20692
rect 16100 20636 16716 20692
rect 16772 20636 21420 20692
rect 21476 20636 21486 20692
rect 28242 20636 28252 20692
rect 28308 20636 29372 20692
rect 29428 20636 29438 20692
rect 29810 20636 29820 20692
rect 29876 20636 30604 20692
rect 30660 20636 33516 20692
rect 33572 20636 34188 20692
rect 34244 20636 34254 20692
rect 35074 20636 35084 20692
rect 35140 20636 36092 20692
rect 36148 20636 36158 20692
rect 41794 20636 41804 20692
rect 41860 20636 44044 20692
rect 44100 20636 47684 20692
rect 52210 20636 52220 20692
rect 52276 20636 55692 20692
rect 55748 20636 56140 20692
rect 56196 20636 56206 20692
rect 29372 20580 29428 20636
rect 7746 20524 7756 20580
rect 7812 20524 10332 20580
rect 10388 20524 10398 20580
rect 22642 20524 22652 20580
rect 22708 20524 25340 20580
rect 25396 20524 25406 20580
rect 29372 20524 31052 20580
rect 31108 20524 31118 20580
rect 42354 20524 42364 20580
rect 42420 20524 44940 20580
rect 44996 20524 47404 20580
rect 47460 20524 47470 20580
rect 47628 20468 47684 20636
rect 47954 20524 47964 20580
rect 48020 20524 53228 20580
rect 53284 20524 53294 20580
rect 6850 20412 6860 20468
rect 6916 20412 9100 20468
rect 9156 20412 10108 20468
rect 10164 20412 10174 20468
rect 16706 20412 16716 20468
rect 16772 20412 21532 20468
rect 21588 20412 21598 20468
rect 47628 20412 48076 20468
rect 48132 20412 52668 20468
rect 52724 20412 52734 20468
rect 15508 20356 15518 20412
rect 15574 20356 15622 20412
rect 15678 20356 15726 20412
rect 15782 20356 15792 20412
rect 29815 20356 29825 20412
rect 29881 20356 29929 20412
rect 29985 20356 30033 20412
rect 30089 20356 30099 20412
rect 44122 20356 44132 20412
rect 44188 20356 44236 20412
rect 44292 20356 44340 20412
rect 44396 20356 44406 20412
rect 58429 20356 58439 20412
rect 58495 20356 58543 20412
rect 58599 20356 58647 20412
rect 58703 20356 58713 20412
rect 2258 20300 2268 20356
rect 2324 20300 2940 20356
rect 2996 20300 3612 20356
rect 3668 20300 5180 20356
rect 5236 20300 5246 20356
rect 30818 20300 30828 20356
rect 30884 20300 34188 20356
rect 34244 20300 34254 20356
rect 59200 20244 60000 20272
rect 2706 20188 2716 20244
rect 2772 20188 2782 20244
rect 8418 20188 8428 20244
rect 8484 20188 10108 20244
rect 10164 20188 11452 20244
rect 11508 20188 11518 20244
rect 18508 20188 20524 20244
rect 20580 20188 20590 20244
rect 26338 20188 26348 20244
rect 26404 20188 29148 20244
rect 29204 20188 29214 20244
rect 30146 20188 30156 20244
rect 30212 20188 36316 20244
rect 36372 20188 37212 20244
rect 37268 20188 37278 20244
rect 42354 20188 42364 20244
rect 42420 20188 43820 20244
rect 43876 20188 44380 20244
rect 44436 20188 45836 20244
rect 45892 20188 45902 20244
rect 50866 20188 50876 20244
rect 50932 20188 52892 20244
rect 52948 20188 53340 20244
rect 53396 20188 53406 20244
rect 57708 20188 60000 20244
rect 2716 20020 2772 20188
rect 18508 20132 18564 20188
rect 57708 20132 57764 20188
rect 59200 20160 60000 20188
rect 9986 20076 9996 20132
rect 10052 20076 15148 20132
rect 15204 20076 15484 20132
rect 15540 20076 15550 20132
rect 15810 20076 15820 20132
rect 15876 20076 16492 20132
rect 16548 20076 16558 20132
rect 16706 20076 16716 20132
rect 16772 20076 18564 20132
rect 26562 20076 26572 20132
rect 26628 20076 38164 20132
rect 38322 20076 38332 20132
rect 38388 20076 38892 20132
rect 38948 20076 38958 20132
rect 45938 20076 45948 20132
rect 46004 20076 47068 20132
rect 47124 20076 47134 20132
rect 47506 20076 47516 20132
rect 47572 20076 50092 20132
rect 50148 20076 50158 20132
rect 54002 20076 54012 20132
rect 54068 20076 55244 20132
rect 55300 20076 55310 20132
rect 57698 20076 57708 20132
rect 57764 20076 57774 20132
rect 38108 20020 38164 20076
rect 2034 19964 2044 20020
rect 2100 19964 3164 20020
rect 3220 19964 3230 20020
rect 3378 19964 3388 20020
rect 3444 19964 4004 20020
rect 7634 19964 7644 20020
rect 7700 19964 10220 20020
rect 10276 19964 10556 20020
rect 10612 19964 11228 20020
rect 11284 19964 11294 20020
rect 12786 19964 12796 20020
rect 12852 19964 15596 20020
rect 15652 19964 15662 20020
rect 17602 19964 17612 20020
rect 17668 19964 21308 20020
rect 21364 19964 21374 20020
rect 24658 19964 24668 20020
rect 24724 19964 25900 20020
rect 25956 19964 25966 20020
rect 30706 19964 30716 20020
rect 30772 19964 33068 20020
rect 33124 19964 33134 20020
rect 36194 19964 36204 20020
rect 36260 19964 37884 20020
rect 37940 19964 37950 20020
rect 38108 19964 39340 20020
rect 39396 19964 39406 20020
rect 40226 19964 40236 20020
rect 40292 19964 42028 20020
rect 42084 19964 42812 20020
rect 42868 19964 42878 20020
rect 46274 19964 46284 20020
rect 46340 19964 46956 20020
rect 47012 19964 47022 20020
rect 49410 19964 49420 20020
rect 49476 19964 52780 20020
rect 52836 19964 52846 20020
rect 2492 19796 2548 19964
rect 3948 19908 4004 19964
rect 3938 19852 3948 19908
rect 4004 19852 4844 19908
rect 4900 19852 4910 19908
rect 7074 19852 7084 19908
rect 7140 19852 8764 19908
rect 8820 19852 8830 19908
rect 9874 19852 9884 19908
rect 9940 19852 19404 19908
rect 19460 19852 19470 19908
rect 20514 19852 20524 19908
rect 20580 19852 21868 19908
rect 21924 19852 21934 19908
rect 35746 19852 35756 19908
rect 35812 19852 38332 19908
rect 38388 19852 38398 19908
rect 38882 19852 38892 19908
rect 38948 19852 40348 19908
rect 40404 19852 40414 19908
rect 42914 19852 42924 19908
rect 42980 19852 43260 19908
rect 43316 19852 43326 19908
rect 47170 19852 47180 19908
rect 47236 19852 49308 19908
rect 49364 19852 49374 19908
rect 2482 19740 2492 19796
rect 2548 19740 2558 19796
rect 29474 19740 29484 19796
rect 29540 19740 35308 19796
rect 35364 19740 35374 19796
rect 35634 19740 35644 19796
rect 35700 19740 37772 19796
rect 37828 19740 42364 19796
rect 42420 19740 42430 19796
rect 45266 19740 45276 19796
rect 45332 19740 46172 19796
rect 46228 19740 51100 19796
rect 51156 19740 52444 19796
rect 52500 19740 52510 19796
rect 15474 19628 15484 19684
rect 15540 19628 17276 19684
rect 17332 19628 17342 19684
rect 46050 19628 46060 19684
rect 46116 19628 46844 19684
rect 46900 19628 48972 19684
rect 49028 19628 49038 19684
rect 8355 19572 8365 19628
rect 8421 19572 8469 19628
rect 8525 19572 8573 19628
rect 8629 19572 8639 19628
rect 22662 19572 22672 19628
rect 22728 19572 22776 19628
rect 22832 19572 22880 19628
rect 22936 19572 22946 19628
rect 36969 19572 36979 19628
rect 37035 19572 37083 19628
rect 37139 19572 37187 19628
rect 37243 19572 37253 19628
rect 51276 19572 51286 19628
rect 51342 19572 51390 19628
rect 51446 19572 51494 19628
rect 51550 19572 51560 19628
rect 16482 19516 16492 19572
rect 16548 19516 21084 19572
rect 21140 19516 21150 19572
rect 23538 19516 23548 19572
rect 23604 19516 23772 19572
rect 23828 19516 25228 19572
rect 25284 19516 25294 19572
rect 46498 19516 46508 19572
rect 46564 19516 47404 19572
rect 47460 19516 47470 19572
rect 8866 19404 8876 19460
rect 8932 19404 10220 19460
rect 10276 19404 10286 19460
rect 15138 19404 15148 19460
rect 15204 19404 16156 19460
rect 16212 19404 16222 19460
rect 17490 19404 17500 19460
rect 17556 19404 17566 19460
rect 24546 19404 24556 19460
rect 24612 19404 26236 19460
rect 26292 19404 26302 19460
rect 34402 19404 34412 19460
rect 34468 19404 34972 19460
rect 35028 19404 36092 19460
rect 36148 19404 36158 19460
rect 43922 19404 43932 19460
rect 43988 19404 46732 19460
rect 46788 19404 46798 19460
rect 0 19348 800 19376
rect 17500 19348 17556 19404
rect 0 19292 1708 19348
rect 1764 19292 4284 19348
rect 4340 19292 4350 19348
rect 16828 19292 17556 19348
rect 26114 19292 26124 19348
rect 26180 19292 27468 19348
rect 27524 19292 27534 19348
rect 30034 19292 30044 19348
rect 30100 19292 33572 19348
rect 51762 19292 51772 19348
rect 51828 19292 53340 19348
rect 53396 19292 54460 19348
rect 54516 19292 54526 19348
rect 0 19264 800 19292
rect 3490 19180 3500 19236
rect 3556 19180 6076 19236
rect 6132 19180 8596 19236
rect 9314 19180 9324 19236
rect 9380 19180 10444 19236
rect 10500 19180 11116 19236
rect 11172 19180 11182 19236
rect 11778 19180 11788 19236
rect 11844 19180 15708 19236
rect 15764 19180 15774 19236
rect 8540 19124 8596 19180
rect 16828 19124 16884 19292
rect 33516 19236 33572 19292
rect 17042 19180 17052 19236
rect 17108 19180 17118 19236
rect 28466 19180 28476 19236
rect 28532 19180 31164 19236
rect 31220 19180 32060 19236
rect 32116 19180 32126 19236
rect 33506 19180 33516 19236
rect 33572 19180 35868 19236
rect 35924 19180 35934 19236
rect 41682 19180 41692 19236
rect 41748 19180 44156 19236
rect 44212 19180 45276 19236
rect 45332 19180 45342 19236
rect 46946 19180 46956 19236
rect 47012 19180 49868 19236
rect 49924 19180 49934 19236
rect 50866 19180 50876 19236
rect 50932 19180 53004 19236
rect 53060 19180 53070 19236
rect 54786 19180 54796 19236
rect 54852 19180 58044 19236
rect 58100 19180 58110 19236
rect 4610 19068 4620 19124
rect 4676 19068 5740 19124
rect 5796 19068 7196 19124
rect 7252 19068 7262 19124
rect 8530 19068 8540 19124
rect 8596 19068 12012 19124
rect 12068 19068 12078 19124
rect 14354 19068 14364 19124
rect 14420 19068 16884 19124
rect 17052 19012 17108 19180
rect 26226 19068 26236 19124
rect 26292 19068 27020 19124
rect 27076 19068 33852 19124
rect 33908 19068 36652 19124
rect 36708 19068 37212 19124
rect 37268 19068 37278 19124
rect 39330 19068 39340 19124
rect 39396 19068 40236 19124
rect 40292 19068 41132 19124
rect 41188 19068 41916 19124
rect 41972 19068 41982 19124
rect 5058 18956 5068 19012
rect 5124 18956 10108 19012
rect 10164 18956 10174 19012
rect 10770 18956 10780 19012
rect 10836 18956 17108 19012
rect 19618 18956 19628 19012
rect 19684 18956 22204 19012
rect 22260 18956 23212 19012
rect 23268 18956 25900 19012
rect 25956 18956 26460 19012
rect 26516 18956 26526 19012
rect 45154 18956 45164 19012
rect 45220 18956 50540 19012
rect 50596 18956 50606 19012
rect 7634 18844 7644 18900
rect 7700 18844 10332 18900
rect 10388 18844 10398 18900
rect 18498 18844 18508 18900
rect 18564 18844 19740 18900
rect 19796 18844 20636 18900
rect 20692 18844 26908 18900
rect 26964 18844 27692 18900
rect 27748 18844 27758 18900
rect 15508 18788 15518 18844
rect 15574 18788 15622 18844
rect 15678 18788 15726 18844
rect 15782 18788 15792 18844
rect 29815 18788 29825 18844
rect 29881 18788 29929 18844
rect 29985 18788 30033 18844
rect 30089 18788 30099 18844
rect 44122 18788 44132 18844
rect 44188 18788 44236 18844
rect 44292 18788 44340 18844
rect 44396 18788 44406 18844
rect 58429 18788 58439 18844
rect 58495 18788 58543 18844
rect 58599 18788 58647 18844
rect 58703 18788 58713 18844
rect 10210 18732 10220 18788
rect 10276 18732 15260 18788
rect 15316 18732 15326 18788
rect 35858 18732 35868 18788
rect 35924 18732 37100 18788
rect 37156 18732 37166 18788
rect 54898 18732 54908 18788
rect 54964 18732 57484 18788
rect 57540 18732 57550 18788
rect 5282 18620 5292 18676
rect 5348 18620 8204 18676
rect 8260 18620 8270 18676
rect 8866 18620 8876 18676
rect 8932 18620 10780 18676
rect 10836 18620 10846 18676
rect 11004 18620 14140 18676
rect 14196 18620 14206 18676
rect 15474 18620 15484 18676
rect 15540 18620 16604 18676
rect 16660 18620 16670 18676
rect 24994 18620 25004 18676
rect 25060 18620 25900 18676
rect 25956 18620 28588 18676
rect 28644 18620 28654 18676
rect 39666 18620 39676 18676
rect 39732 18620 40460 18676
rect 40516 18620 41468 18676
rect 41524 18620 41534 18676
rect 48860 18620 49756 18676
rect 49812 18620 49822 18676
rect 11004 18564 11060 18620
rect 48860 18564 48916 18620
rect 3938 18508 3948 18564
rect 4004 18508 5740 18564
rect 5796 18508 6748 18564
rect 6804 18508 6814 18564
rect 7074 18508 7084 18564
rect 7140 18508 7420 18564
rect 7476 18508 7486 18564
rect 9090 18508 9100 18564
rect 9156 18508 9166 18564
rect 10322 18508 10332 18564
rect 10388 18508 11060 18564
rect 12450 18508 12460 18564
rect 12516 18508 14700 18564
rect 14756 18508 14766 18564
rect 15250 18508 15260 18564
rect 15316 18508 16492 18564
rect 16548 18508 16558 18564
rect 18274 18508 18284 18564
rect 18340 18508 19292 18564
rect 19348 18508 19358 18564
rect 22082 18508 22092 18564
rect 22148 18508 22540 18564
rect 22596 18508 23436 18564
rect 23492 18508 23502 18564
rect 26562 18508 26572 18564
rect 26628 18508 28700 18564
rect 28756 18508 29708 18564
rect 29764 18508 29774 18564
rect 31938 18508 31948 18564
rect 32004 18508 34748 18564
rect 34804 18508 34814 18564
rect 41234 18508 41244 18564
rect 41300 18508 42812 18564
rect 42868 18508 42878 18564
rect 48178 18508 48188 18564
rect 48244 18508 48860 18564
rect 48916 18508 48926 18564
rect 49410 18508 49420 18564
rect 49476 18508 52332 18564
rect 52388 18508 52398 18564
rect 54450 18508 54460 18564
rect 54516 18508 55132 18564
rect 55188 18508 55198 18564
rect 9100 18452 9156 18508
rect 2818 18396 2828 18452
rect 2884 18396 3836 18452
rect 3892 18396 4396 18452
rect 4452 18396 4462 18452
rect 6066 18396 6076 18452
rect 6132 18396 6972 18452
rect 7028 18396 7038 18452
rect 9100 18396 13692 18452
rect 13748 18396 13758 18452
rect 15092 18396 16828 18452
rect 16884 18396 17388 18452
rect 17444 18396 17454 18452
rect 18834 18396 18844 18452
rect 18900 18396 20748 18452
rect 20804 18396 21308 18452
rect 21364 18396 21374 18452
rect 24210 18396 24220 18452
rect 24276 18396 25228 18452
rect 25284 18396 25294 18452
rect 27346 18396 27356 18452
rect 27412 18396 29148 18452
rect 29204 18396 29214 18452
rect 33394 18396 33404 18452
rect 33460 18396 35196 18452
rect 35252 18396 35756 18452
rect 35812 18396 35822 18452
rect 36082 18396 36092 18452
rect 36148 18396 37100 18452
rect 37156 18396 37166 18452
rect 38612 18396 38780 18452
rect 38836 18396 38846 18452
rect 42914 18396 42924 18452
rect 42980 18396 46732 18452
rect 46788 18396 47628 18452
rect 47684 18396 47694 18452
rect 48066 18396 48076 18452
rect 48132 18396 52556 18452
rect 52612 18396 52622 18452
rect 6076 18340 6132 18396
rect 15092 18340 15148 18396
rect 38612 18340 38668 18396
rect 1922 18284 1932 18340
rect 1988 18284 6132 18340
rect 7074 18284 7084 18340
rect 7140 18284 9660 18340
rect 9716 18284 9726 18340
rect 10994 18284 11004 18340
rect 11060 18284 11564 18340
rect 11620 18284 11630 18340
rect 12002 18284 12012 18340
rect 12068 18284 15148 18340
rect 16930 18284 16940 18340
rect 16996 18284 17724 18340
rect 17780 18284 17790 18340
rect 18722 18284 18732 18340
rect 18788 18284 22764 18340
rect 22820 18284 23324 18340
rect 23380 18284 23390 18340
rect 24658 18284 24668 18340
rect 24724 18284 25564 18340
rect 25620 18284 25630 18340
rect 27346 18284 27356 18340
rect 27412 18284 27916 18340
rect 27972 18284 27982 18340
rect 35074 18284 35084 18340
rect 35140 18284 35868 18340
rect 35924 18284 35934 18340
rect 36530 18284 36540 18340
rect 36596 18284 38668 18340
rect 40338 18284 40348 18340
rect 40404 18284 41524 18340
rect 41794 18284 41804 18340
rect 41860 18284 44604 18340
rect 44660 18284 46844 18340
rect 46900 18284 46910 18340
rect 49186 18284 49196 18340
rect 49252 18284 49532 18340
rect 49588 18284 49598 18340
rect 53890 18284 53900 18340
rect 53956 18284 54236 18340
rect 54292 18284 54302 18340
rect 41468 18228 41524 18284
rect 7970 18172 7980 18228
rect 8036 18172 10500 18228
rect 10658 18172 10668 18228
rect 10724 18172 12348 18228
rect 12404 18172 12414 18228
rect 15810 18172 15820 18228
rect 15876 18172 16156 18228
rect 16212 18172 16222 18228
rect 26852 18172 40404 18228
rect 41468 18172 42140 18228
rect 42196 18172 48748 18228
rect 48804 18172 48814 18228
rect 10444 18116 10500 18172
rect 10444 18060 11228 18116
rect 11284 18060 11294 18116
rect 8355 18004 8365 18060
rect 8421 18004 8469 18060
rect 8525 18004 8573 18060
rect 8629 18004 8639 18060
rect 22662 18004 22672 18060
rect 22728 18004 22776 18060
rect 22832 18004 22880 18060
rect 22936 18004 22946 18060
rect 26852 18004 26908 18172
rect 34514 18060 34524 18116
rect 34580 18060 34860 18116
rect 34916 18060 34926 18116
rect 36969 18004 36979 18060
rect 37035 18004 37083 18060
rect 37139 18004 37187 18060
rect 37243 18004 37253 18060
rect 25330 17948 25340 18004
rect 25396 17948 26908 18004
rect 7186 17836 7196 17892
rect 7252 17836 8204 17892
rect 8260 17836 11900 17892
rect 11956 17836 11966 17892
rect 15026 17836 15036 17892
rect 15092 17836 20412 17892
rect 20468 17836 21868 17892
rect 21924 17836 23100 17892
rect 23156 17836 23166 17892
rect 27906 17836 27916 17892
rect 27972 17836 28028 17892
rect 28084 17836 28094 17892
rect 37548 17836 39564 17892
rect 39620 17836 39630 17892
rect 2034 17724 2044 17780
rect 2100 17724 2940 17780
rect 2996 17724 3612 17780
rect 3668 17724 5628 17780
rect 5684 17724 5694 17780
rect 6066 17724 6076 17780
rect 6132 17724 7084 17780
rect 7140 17724 7150 17780
rect 7970 17724 7980 17780
rect 8036 17724 11004 17780
rect 11060 17724 11070 17780
rect 12012 17724 17500 17780
rect 17556 17724 17566 17780
rect 26450 17724 26460 17780
rect 26516 17724 28420 17780
rect 8306 17612 8316 17668
rect 8372 17612 11788 17668
rect 11844 17612 11854 17668
rect 0 17556 800 17584
rect 12012 17556 12068 17724
rect 28364 17668 28420 17724
rect 37548 17668 37604 17836
rect 40348 17780 40404 18172
rect 49196 18116 49252 18284
rect 41234 18060 41244 18116
rect 41300 18060 41580 18116
rect 41636 18060 41646 18116
rect 43250 18060 43260 18116
rect 43316 18060 45276 18116
rect 45332 18060 49252 18116
rect 51276 18004 51286 18060
rect 51342 18004 51390 18060
rect 51446 18004 51494 18060
rect 51550 18004 51560 18060
rect 42242 17836 42252 17892
rect 42308 17836 42812 17892
rect 42868 17836 42878 17892
rect 53218 17836 53228 17892
rect 53284 17836 54012 17892
rect 54068 17836 54572 17892
rect 54628 17836 54638 17892
rect 38612 17724 39004 17780
rect 39060 17724 39070 17780
rect 40338 17724 40348 17780
rect 40404 17724 41020 17780
rect 41076 17724 41692 17780
rect 41748 17724 41758 17780
rect 53106 17724 53116 17780
rect 53172 17724 53564 17780
rect 53620 17724 53630 17780
rect 12898 17612 12908 17668
rect 12964 17612 18172 17668
rect 18228 17612 18238 17668
rect 21522 17612 21532 17668
rect 21588 17612 28196 17668
rect 28354 17612 28364 17668
rect 28420 17612 30380 17668
rect 30436 17612 30446 17668
rect 31154 17612 31164 17668
rect 31220 17612 37548 17668
rect 37604 17612 37614 17668
rect 0 17500 1820 17556
rect 1876 17500 1886 17556
rect 10098 17500 10108 17556
rect 10164 17500 12068 17556
rect 18172 17556 18228 17612
rect 28140 17556 28196 17612
rect 38612 17556 38668 17724
rect 44706 17612 44716 17668
rect 44772 17612 46284 17668
rect 46340 17612 46350 17668
rect 18172 17500 21420 17556
rect 21476 17500 21486 17556
rect 23202 17500 23212 17556
rect 23268 17500 24332 17556
rect 24388 17500 24398 17556
rect 26002 17500 26012 17556
rect 26068 17500 27692 17556
rect 27748 17500 27758 17556
rect 28140 17500 34524 17556
rect 34580 17500 35756 17556
rect 35812 17500 37100 17556
rect 37156 17500 38668 17556
rect 0 17472 800 17500
rect 4498 17388 4508 17444
rect 4564 17388 4732 17444
rect 4788 17388 5516 17444
rect 5572 17388 5582 17444
rect 10434 17388 10444 17444
rect 10500 17388 11676 17444
rect 11732 17388 18396 17444
rect 18452 17388 18462 17444
rect 25330 17388 25340 17444
rect 25396 17388 26236 17444
rect 26292 17388 26302 17444
rect 35522 17388 35532 17444
rect 35588 17388 37548 17444
rect 37604 17388 37614 17444
rect 42242 17388 42252 17444
rect 42308 17388 43148 17444
rect 43204 17388 43214 17444
rect 51650 17388 51660 17444
rect 51716 17388 51996 17444
rect 52052 17388 54068 17444
rect 54226 17388 54236 17444
rect 54292 17388 55244 17444
rect 55300 17388 57036 17444
rect 57092 17388 57102 17444
rect 54012 17332 54068 17388
rect 8082 17276 8092 17332
rect 8148 17276 9772 17332
rect 9828 17276 9838 17332
rect 12338 17276 12348 17332
rect 12404 17276 15148 17332
rect 19394 17276 19404 17332
rect 19460 17276 27356 17332
rect 27412 17276 27422 17332
rect 42466 17276 42476 17332
rect 42532 17276 42542 17332
rect 54012 17276 54796 17332
rect 54852 17276 55356 17332
rect 55412 17276 55422 17332
rect 2258 17052 2268 17108
rect 2324 17052 3052 17108
rect 3108 17052 3118 17108
rect 3332 16884 3388 17220
rect 3444 17164 3454 17220
rect 13010 17164 13020 17220
rect 13076 17164 14364 17220
rect 14420 17164 14430 17220
rect 7074 17052 7084 17108
rect 7140 17052 9100 17108
rect 9156 17052 9166 17108
rect 12898 17052 12908 17108
rect 12964 17052 14588 17108
rect 14644 17052 14654 17108
rect 15092 16996 15148 17276
rect 15508 17220 15518 17276
rect 15574 17220 15622 17276
rect 15678 17220 15726 17276
rect 15782 17220 15792 17276
rect 29815 17220 29825 17276
rect 29881 17220 29929 17276
rect 29985 17220 30033 17276
rect 30089 17220 30099 17276
rect 23538 17164 23548 17220
rect 23604 17164 28364 17220
rect 28420 17164 28430 17220
rect 33058 17164 33068 17220
rect 33124 17164 33740 17220
rect 33796 17164 36316 17220
rect 36372 17164 36382 17220
rect 42476 17108 42532 17276
rect 44122 17220 44132 17276
rect 44188 17220 44236 17276
rect 44292 17220 44340 17276
rect 44396 17220 44406 17276
rect 58429 17220 58439 17276
rect 58495 17220 58543 17276
rect 58599 17220 58647 17276
rect 58703 17220 58713 17276
rect 23324 17052 23772 17108
rect 23828 17052 23838 17108
rect 24434 17052 24444 17108
rect 24500 17052 26460 17108
rect 26516 17052 26526 17108
rect 32050 17052 32060 17108
rect 32116 17052 33516 17108
rect 33572 17052 33582 17108
rect 34290 17052 34300 17108
rect 34356 17052 34972 17108
rect 35028 17052 35038 17108
rect 40450 17052 40460 17108
rect 40516 17052 41244 17108
rect 41300 17052 41310 17108
rect 42130 17052 42140 17108
rect 42196 17052 45388 17108
rect 45444 17052 49308 17108
rect 49364 17052 49374 17108
rect 53554 17052 53564 17108
rect 53620 17052 58156 17108
rect 58212 17052 58222 17108
rect 23324 16996 23380 17052
rect 4610 16940 4620 16996
rect 4676 16940 5740 16996
rect 5796 16940 7140 16996
rect 7858 16940 7868 16996
rect 7924 16940 9044 16996
rect 10994 16940 11004 16996
rect 11060 16940 13412 16996
rect 15092 16940 15596 16996
rect 15652 16940 15662 16996
rect 22418 16940 22428 16996
rect 22484 16940 23324 16996
rect 23380 16940 23390 16996
rect 25554 16940 25564 16996
rect 25620 16940 27244 16996
rect 27300 16940 29260 16996
rect 29316 16940 33068 16996
rect 33124 16940 33134 16996
rect 7084 16884 7140 16940
rect 8988 16884 9044 16940
rect 2258 16828 2268 16884
rect 2324 16828 3388 16884
rect 3714 16828 3724 16884
rect 3780 16828 4508 16884
rect 4564 16828 6524 16884
rect 6580 16828 6590 16884
rect 7074 16828 7084 16884
rect 7140 16828 8764 16884
rect 8820 16828 8830 16884
rect 8978 16828 8988 16884
rect 9044 16828 9660 16884
rect 9716 16828 9726 16884
rect 2034 16716 2044 16772
rect 2100 16716 2940 16772
rect 2996 16716 3500 16772
rect 3556 16716 3566 16772
rect 5282 16716 5292 16772
rect 5348 16716 6076 16772
rect 6132 16716 6142 16772
rect 7858 16716 7868 16772
rect 7924 16716 9772 16772
rect 9828 16716 10892 16772
rect 10948 16716 10958 16772
rect 13356 16548 13412 16940
rect 33516 16884 33572 17052
rect 42588 16884 42644 17052
rect 50978 16940 50988 16996
rect 51044 16940 52108 16996
rect 52164 16940 53900 16996
rect 53956 16940 53966 16996
rect 18722 16828 18732 16884
rect 18788 16828 19292 16884
rect 19348 16828 19358 16884
rect 19506 16828 19516 16884
rect 19572 16828 20412 16884
rect 20468 16828 20478 16884
rect 26338 16828 26348 16884
rect 26404 16828 27692 16884
rect 27748 16828 27758 16884
rect 29586 16828 29596 16884
rect 29652 16828 32172 16884
rect 32228 16828 33292 16884
rect 33348 16828 33358 16884
rect 33516 16828 34636 16884
rect 34692 16828 34702 16884
rect 41570 16828 41580 16884
rect 41636 16828 41646 16884
rect 42578 16828 42588 16884
rect 42644 16828 42654 16884
rect 56466 16828 56476 16884
rect 56532 16828 57932 16884
rect 57988 16828 57998 16884
rect 41580 16772 41636 16828
rect 19730 16716 19740 16772
rect 19796 16716 23212 16772
rect 23268 16716 23278 16772
rect 30706 16716 30716 16772
rect 30772 16716 31724 16772
rect 31780 16716 31790 16772
rect 32732 16716 39228 16772
rect 39284 16716 39294 16772
rect 41580 16716 43708 16772
rect 43764 16716 43774 16772
rect 50418 16716 50428 16772
rect 50484 16716 51548 16772
rect 51604 16716 51614 16772
rect 51762 16716 51772 16772
rect 51828 16716 53340 16772
rect 53396 16716 53406 16772
rect 53890 16716 53900 16772
rect 53956 16716 55580 16772
rect 55636 16716 56924 16772
rect 56980 16716 56990 16772
rect 32732 16660 32788 16716
rect 59200 16660 60000 16688
rect 16594 16604 16604 16660
rect 16660 16604 17164 16660
rect 17220 16604 17230 16660
rect 24322 16604 24332 16660
rect 24388 16604 32788 16660
rect 33506 16604 33516 16660
rect 33572 16604 33852 16660
rect 33908 16604 33918 16660
rect 36754 16604 36764 16660
rect 36820 16604 37772 16660
rect 37828 16604 37838 16660
rect 57138 16604 57148 16660
rect 57204 16604 57596 16660
rect 57652 16604 57662 16660
rect 58034 16604 58044 16660
rect 58100 16604 60000 16660
rect 33516 16548 33572 16604
rect 59200 16576 60000 16604
rect 2706 16492 2716 16548
rect 2772 16492 5292 16548
rect 5348 16492 5358 16548
rect 13356 16492 20748 16548
rect 20804 16492 20814 16548
rect 24770 16492 24780 16548
rect 24836 16492 27916 16548
rect 27972 16492 28252 16548
rect 28308 16492 28318 16548
rect 30258 16492 30268 16548
rect 30324 16492 31500 16548
rect 31556 16492 33572 16548
rect 8355 16436 8365 16492
rect 8421 16436 8469 16492
rect 8525 16436 8573 16492
rect 8629 16436 8639 16492
rect 22662 16436 22672 16492
rect 22728 16436 22776 16492
rect 22832 16436 22880 16492
rect 22936 16436 22946 16492
rect 36969 16436 36979 16492
rect 37035 16436 37083 16492
rect 37139 16436 37187 16492
rect 37243 16436 37253 16492
rect 51276 16436 51286 16492
rect 51342 16436 51390 16492
rect 51446 16436 51494 16492
rect 51550 16436 51560 16492
rect 2258 16380 2268 16436
rect 2324 16380 3164 16436
rect 3220 16380 3230 16436
rect 10882 16380 10892 16436
rect 10948 16380 13468 16436
rect 13524 16380 13534 16436
rect 26114 16380 26124 16436
rect 26180 16380 27020 16436
rect 27076 16380 29596 16436
rect 29652 16380 29662 16436
rect 55010 16380 55020 16436
rect 55076 16380 55468 16436
rect 55524 16380 55534 16436
rect 2482 16268 2492 16324
rect 2548 16268 6132 16324
rect 9986 16268 9996 16324
rect 10052 16268 20412 16324
rect 20468 16268 20478 16324
rect 54562 16268 54572 16324
rect 54628 16268 55692 16324
rect 55748 16268 55758 16324
rect 6076 16212 6132 16268
rect 3378 16156 3388 16212
rect 3444 16156 4172 16212
rect 4228 16156 4238 16212
rect 6066 16156 6076 16212
rect 6132 16156 6524 16212
rect 6580 16156 6590 16212
rect 8082 16156 8092 16212
rect 8148 16156 21084 16212
rect 21140 16156 21150 16212
rect 23426 16156 23436 16212
rect 23492 16156 33740 16212
rect 33796 16156 34860 16212
rect 34916 16156 34926 16212
rect 36418 16156 36428 16212
rect 36484 16156 38836 16212
rect 51426 16156 51436 16212
rect 51492 16156 53228 16212
rect 53284 16156 53676 16212
rect 53732 16156 53742 16212
rect 54674 16156 54684 16212
rect 54740 16156 55580 16212
rect 55636 16156 55646 16212
rect 6524 16100 6580 16156
rect 38780 16100 38836 16156
rect 6524 16044 8540 16100
rect 8596 16044 8606 16100
rect 12338 16044 12348 16100
rect 12404 16044 13356 16100
rect 13412 16044 13422 16100
rect 18834 16044 18844 16100
rect 18900 16044 20076 16100
rect 20132 16044 20142 16100
rect 21522 16044 21532 16100
rect 21588 16044 22204 16100
rect 22260 16044 22270 16100
rect 23202 16044 23212 16100
rect 23268 16044 23884 16100
rect 23940 16044 24556 16100
rect 24612 16044 25452 16100
rect 25508 16044 25518 16100
rect 27122 16044 27132 16100
rect 27188 16044 27356 16100
rect 27412 16044 28140 16100
rect 28196 16044 28206 16100
rect 36978 16044 36988 16100
rect 37044 16044 37884 16100
rect 37940 16044 37950 16100
rect 38770 16044 38780 16100
rect 38836 16044 38846 16100
rect 43922 16044 43932 16100
rect 43988 16044 45052 16100
rect 45108 16044 45118 16100
rect 48962 16044 48972 16100
rect 49028 16044 51660 16100
rect 51716 16044 51884 16100
rect 51940 16044 51950 16100
rect 54338 16044 54348 16100
rect 54404 16044 54908 16100
rect 54964 16044 54974 16100
rect 55346 16044 55356 16100
rect 55412 16044 57372 16100
rect 57428 16044 57438 16100
rect 13570 15932 13580 15988
rect 13636 15932 14476 15988
rect 14532 15932 18060 15988
rect 18116 15932 18126 15988
rect 20076 15876 20132 16044
rect 55356 15988 55412 16044
rect 20962 15932 20972 15988
rect 21028 15932 21980 15988
rect 22036 15932 22046 15988
rect 28578 15932 28588 15988
rect 28644 15932 35084 15988
rect 35140 15932 36092 15988
rect 36148 15932 36158 15988
rect 45826 15932 45836 15988
rect 45892 15932 46508 15988
rect 46564 15932 47628 15988
rect 47684 15932 47964 15988
rect 48020 15932 49308 15988
rect 49364 15932 51772 15988
rect 51828 15932 51838 15988
rect 55010 15932 55020 15988
rect 55076 15932 55412 15988
rect 13906 15820 13916 15876
rect 13972 15820 15036 15876
rect 15092 15820 15102 15876
rect 20076 15820 22316 15876
rect 22372 15820 22382 15876
rect 24546 15820 24556 15876
rect 24612 15820 26012 15876
rect 26068 15820 26684 15876
rect 26740 15820 26750 15876
rect 28466 15820 28476 15876
rect 28532 15820 32060 15876
rect 32116 15820 32126 15876
rect 43810 15820 43820 15876
rect 43876 15820 45724 15876
rect 45780 15820 45790 15876
rect 50418 15820 50428 15876
rect 50484 15820 50652 15876
rect 50708 15820 50718 15876
rect 0 15764 800 15792
rect 0 15708 1596 15764
rect 1652 15708 1662 15764
rect 26898 15708 26908 15764
rect 26964 15708 27692 15764
rect 27748 15708 28364 15764
rect 28420 15708 28430 15764
rect 0 15680 800 15708
rect 15508 15652 15518 15708
rect 15574 15652 15622 15708
rect 15678 15652 15726 15708
rect 15782 15652 15792 15708
rect 29815 15652 29825 15708
rect 29881 15652 29929 15708
rect 29985 15652 30033 15708
rect 30089 15652 30099 15708
rect 44122 15652 44132 15708
rect 44188 15652 44236 15708
rect 44292 15652 44340 15708
rect 44396 15652 44406 15708
rect 58429 15652 58439 15708
rect 58495 15652 58543 15708
rect 58599 15652 58647 15708
rect 58703 15652 58713 15708
rect 7410 15596 7420 15652
rect 7476 15596 10556 15652
rect 10612 15596 11004 15652
rect 11060 15596 11070 15652
rect 4722 15484 4732 15540
rect 4788 15484 26908 15540
rect 27010 15484 27020 15540
rect 27076 15484 30268 15540
rect 30324 15484 30334 15540
rect 34178 15484 34188 15540
rect 34244 15484 35196 15540
rect 35252 15484 35262 15540
rect 40226 15484 40236 15540
rect 40292 15484 42140 15540
rect 42196 15484 42206 15540
rect 44594 15484 44604 15540
rect 44660 15484 45388 15540
rect 45444 15484 50428 15540
rect 50484 15484 50494 15540
rect 54786 15484 54796 15540
rect 54852 15484 55244 15540
rect 55300 15484 55310 15540
rect 26852 15428 26908 15484
rect 2258 15372 2268 15428
rect 2324 15372 2604 15428
rect 2660 15372 2828 15428
rect 2884 15372 2894 15428
rect 3332 15372 3500 15428
rect 3556 15372 4396 15428
rect 4452 15372 4462 15428
rect 5282 15372 5292 15428
rect 5348 15372 6636 15428
rect 6692 15372 6702 15428
rect 6860 15372 7084 15428
rect 7140 15372 8988 15428
rect 9044 15372 9660 15428
rect 9716 15372 9726 15428
rect 12002 15372 12012 15428
rect 12068 15372 15148 15428
rect 15204 15372 15484 15428
rect 15540 15372 16268 15428
rect 16324 15372 16334 15428
rect 26852 15372 47068 15428
rect 47842 15372 47852 15428
rect 47908 15372 51436 15428
rect 51492 15372 51502 15428
rect 1922 15260 1932 15316
rect 1988 15260 2716 15316
rect 2772 15260 2782 15316
rect 3332 15204 3388 15372
rect 2604 15148 3388 15204
rect 2604 15092 2660 15148
rect 6860 15092 6916 15372
rect 47012 15316 47068 15372
rect 11666 15260 11676 15316
rect 11732 15260 12348 15316
rect 12404 15260 12414 15316
rect 12674 15260 12684 15316
rect 12740 15260 14140 15316
rect 14196 15260 14206 15316
rect 14914 15260 14924 15316
rect 14980 15260 16380 15316
rect 16436 15260 16446 15316
rect 28242 15260 28252 15316
rect 28308 15260 30828 15316
rect 30884 15260 30894 15316
rect 33954 15260 33964 15316
rect 34020 15260 34972 15316
rect 35028 15260 35038 15316
rect 37314 15260 37324 15316
rect 37380 15260 40908 15316
rect 40964 15260 40974 15316
rect 41234 15260 41244 15316
rect 41300 15260 41580 15316
rect 41636 15260 42364 15316
rect 42420 15260 42430 15316
rect 47012 15260 47516 15316
rect 47572 15260 50652 15316
rect 50708 15260 50718 15316
rect 51202 15260 51212 15316
rect 51268 15260 51772 15316
rect 51828 15260 51838 15316
rect 53442 15260 53452 15316
rect 53508 15260 55132 15316
rect 55188 15260 55198 15316
rect 16146 15148 16156 15204
rect 16212 15148 17724 15204
rect 17780 15148 17790 15204
rect 22418 15148 22428 15204
rect 22484 15148 24108 15204
rect 24164 15148 24174 15204
rect 31714 15148 31724 15204
rect 31780 15148 36988 15204
rect 37044 15148 37054 15204
rect 39330 15148 39340 15204
rect 39396 15148 40012 15204
rect 40068 15148 40078 15204
rect 48178 15148 48188 15204
rect 48244 15148 49196 15204
rect 49252 15148 49262 15204
rect 50418 15148 50428 15204
rect 50484 15148 50522 15204
rect 53778 15148 53788 15204
rect 53844 15148 54012 15204
rect 54068 15148 54078 15204
rect 2594 15036 2604 15092
rect 2660 15036 2670 15092
rect 5954 15036 5964 15092
rect 6020 15036 6916 15092
rect 7084 15036 23492 15092
rect 35858 15036 35868 15092
rect 35924 15036 37100 15092
rect 37156 15036 37166 15092
rect 49858 15036 49868 15092
rect 49924 15036 50092 15092
rect 50148 15036 50158 15092
rect 7084 14980 7140 15036
rect 23436 14980 23492 15036
rect 4498 14924 4508 14980
rect 4564 14924 5516 14980
rect 5572 14924 6300 14980
rect 6356 14924 7140 14980
rect 23426 14924 23436 14980
rect 23492 14924 24780 14980
rect 24836 14924 24846 14980
rect 32498 14924 32508 14980
rect 32564 14924 33516 14980
rect 33572 14924 35756 14980
rect 35812 14924 35822 14980
rect 53890 14924 53900 14980
rect 53956 14924 54572 14980
rect 54628 14924 54638 14980
rect 8355 14868 8365 14924
rect 8421 14868 8469 14924
rect 8525 14868 8573 14924
rect 8629 14868 8639 14924
rect 22662 14868 22672 14924
rect 22728 14868 22776 14924
rect 22832 14868 22880 14924
rect 22936 14868 22946 14924
rect 36969 14868 36979 14924
rect 37035 14868 37083 14924
rect 37139 14868 37187 14924
rect 37243 14868 37253 14924
rect 51276 14868 51286 14924
rect 51342 14868 51390 14924
rect 51446 14868 51494 14924
rect 51550 14868 51560 14924
rect 1810 14812 1820 14868
rect 1876 14812 1886 14868
rect 2146 14812 2156 14868
rect 2212 14812 3164 14868
rect 3220 14812 3230 14868
rect 9986 14812 9996 14868
rect 10052 14812 11452 14868
rect 11508 14812 14252 14868
rect 14308 14812 16940 14868
rect 16996 14812 18172 14868
rect 18228 14812 18620 14868
rect 18676 14812 18686 14868
rect 18946 14812 18956 14868
rect 19012 14812 20300 14868
rect 20356 14812 20366 14868
rect 53442 14812 53452 14868
rect 53508 14812 55132 14868
rect 55188 14812 56252 14868
rect 56308 14812 56318 14868
rect 1820 14644 1876 14812
rect 8978 14700 8988 14756
rect 9044 14700 9884 14756
rect 9940 14700 9950 14756
rect 26786 14700 26796 14756
rect 26852 14700 42700 14756
rect 42756 14700 42766 14756
rect 50418 14700 50428 14756
rect 50484 14700 51884 14756
rect 51940 14700 51950 14756
rect 1810 14588 1820 14644
rect 1876 14588 1886 14644
rect 10994 14588 11004 14644
rect 11060 14588 13468 14644
rect 13524 14588 13804 14644
rect 13860 14588 19404 14644
rect 19460 14588 19470 14644
rect 21522 14588 21532 14644
rect 21588 14588 23884 14644
rect 23940 14588 25116 14644
rect 25172 14588 25182 14644
rect 28466 14588 28476 14644
rect 28532 14588 38668 14644
rect 39554 14588 39564 14644
rect 39620 14588 40572 14644
rect 40628 14588 40638 14644
rect 38612 14532 38668 14588
rect 2930 14476 2940 14532
rect 2996 14476 4284 14532
rect 4340 14476 4350 14532
rect 6178 14476 6188 14532
rect 6244 14476 6636 14532
rect 6692 14476 6702 14532
rect 11442 14476 11452 14532
rect 11508 14476 12124 14532
rect 12180 14476 12190 14532
rect 15250 14476 15260 14532
rect 15316 14476 16044 14532
rect 16100 14476 16110 14532
rect 19618 14476 19628 14532
rect 19684 14476 21868 14532
rect 21924 14476 23324 14532
rect 23380 14476 23390 14532
rect 23538 14476 23548 14532
rect 23604 14476 24444 14532
rect 24500 14476 24510 14532
rect 27458 14476 27468 14532
rect 27524 14476 28252 14532
rect 28308 14476 28318 14532
rect 31154 14476 31164 14532
rect 31220 14476 32396 14532
rect 32452 14476 32462 14532
rect 36978 14476 36988 14532
rect 37044 14476 37884 14532
rect 37940 14476 37950 14532
rect 38612 14476 44268 14532
rect 44324 14476 44828 14532
rect 44884 14476 44894 14532
rect 55794 14476 55804 14532
rect 55860 14476 56476 14532
rect 56532 14476 57260 14532
rect 57316 14476 57326 14532
rect 6188 14420 6244 14476
rect 3938 14364 3948 14420
rect 4004 14364 6244 14420
rect 6402 14364 6412 14420
rect 6468 14364 10332 14420
rect 10388 14364 11564 14420
rect 11620 14364 14252 14420
rect 14308 14364 16604 14420
rect 16660 14364 16670 14420
rect 17154 14364 17164 14420
rect 17220 14364 18396 14420
rect 18452 14364 18462 14420
rect 34402 14364 34412 14420
rect 34468 14364 35868 14420
rect 35924 14364 35934 14420
rect 38322 14364 38332 14420
rect 38388 14364 39228 14420
rect 39284 14364 39900 14420
rect 39956 14364 39966 14420
rect 44594 14364 44604 14420
rect 44660 14364 45276 14420
rect 45332 14364 45342 14420
rect 45826 14364 45836 14420
rect 45892 14364 47516 14420
rect 47572 14364 47582 14420
rect 55346 14364 55356 14420
rect 55412 14364 57036 14420
rect 57092 14364 57102 14420
rect 6738 14252 6748 14308
rect 6804 14252 8204 14308
rect 8260 14252 9436 14308
rect 9492 14252 9502 14308
rect 16034 14252 16044 14308
rect 16100 14252 16716 14308
rect 16772 14252 16782 14308
rect 36194 14252 36204 14308
rect 36260 14252 50540 14308
rect 50596 14252 50606 14308
rect 52098 14252 52108 14308
rect 52164 14252 53004 14308
rect 53060 14252 53788 14308
rect 53844 14252 53854 14308
rect 54562 14252 54572 14308
rect 54628 14252 54638 14308
rect 54572 14196 54628 14252
rect 3602 14140 3612 14196
rect 3668 14140 4172 14196
rect 4228 14140 4238 14196
rect 5618 14140 5628 14196
rect 5684 14140 9772 14196
rect 9828 14140 9838 14196
rect 16268 14140 22988 14196
rect 23044 14140 23772 14196
rect 23828 14140 23838 14196
rect 25900 14140 26796 14196
rect 26852 14140 26862 14196
rect 37538 14140 37548 14196
rect 37604 14140 38220 14196
rect 38276 14140 38286 14196
rect 38658 14140 38668 14196
rect 38724 14140 39452 14196
rect 39508 14140 39518 14196
rect 48178 14140 48188 14196
rect 48244 14140 48748 14196
rect 48804 14140 54628 14196
rect 15508 14084 15518 14140
rect 15574 14084 15622 14140
rect 15678 14084 15726 14140
rect 15782 14084 15792 14140
rect 2258 14028 2268 14084
rect 2324 14028 8036 14084
rect 0 13972 800 14000
rect 0 13916 1708 13972
rect 1764 13916 1774 13972
rect 4274 13916 4284 13972
rect 4340 13916 6860 13972
rect 6916 13916 6926 13972
rect 0 13888 800 13916
rect 2706 13804 2716 13860
rect 2772 13804 5964 13860
rect 6020 13804 6030 13860
rect 7980 13748 8036 14028
rect 15698 13916 15708 13972
rect 15764 13916 16044 13972
rect 16100 13916 16110 13972
rect 10770 13804 10780 13860
rect 10836 13804 14812 13860
rect 14868 13804 14878 13860
rect 15026 13804 15036 13860
rect 15092 13804 15596 13860
rect 15652 13804 15662 13860
rect 16268 13748 16324 14140
rect 16594 14028 16604 14084
rect 16660 14028 16940 14084
rect 16996 14028 17006 14084
rect 25900 13972 25956 14140
rect 29815 14084 29825 14140
rect 29881 14084 29929 14140
rect 29985 14084 30033 14140
rect 30089 14084 30099 14140
rect 44122 14084 44132 14140
rect 44188 14084 44236 14140
rect 44292 14084 44340 14140
rect 44396 14084 44406 14140
rect 58429 14084 58439 14140
rect 58495 14084 58543 14140
rect 58599 14084 58647 14140
rect 58703 14084 58713 14140
rect 49410 14028 49420 14084
rect 49476 14028 49868 14084
rect 49924 14028 53228 14084
rect 53284 14028 55244 14084
rect 55300 14028 56140 14084
rect 56196 14028 56206 14084
rect 16482 13916 16492 13972
rect 16548 13916 17388 13972
rect 17444 13916 17454 13972
rect 18274 13916 18284 13972
rect 18340 13916 19068 13972
rect 19124 13916 19134 13972
rect 24770 13916 24780 13972
rect 24836 13916 25900 13972
rect 25956 13916 25966 13972
rect 27122 13916 27132 13972
rect 27188 13916 27692 13972
rect 27748 13916 27758 13972
rect 41234 13916 41244 13972
rect 41300 13916 41692 13972
rect 41748 13916 41758 13972
rect 55878 13916 55916 13972
rect 55972 13916 55982 13972
rect 16594 13804 16604 13860
rect 16660 13804 16716 13860
rect 16772 13804 17612 13860
rect 17668 13804 17678 13860
rect 18386 13804 18396 13860
rect 18452 13804 21196 13860
rect 21252 13804 21644 13860
rect 21700 13804 23100 13860
rect 23156 13804 23166 13860
rect 28578 13804 28588 13860
rect 28644 13804 30044 13860
rect 30100 13804 30110 13860
rect 36082 13804 36092 13860
rect 36148 13804 37884 13860
rect 37940 13804 37950 13860
rect 39554 13804 39564 13860
rect 39620 13804 41580 13860
rect 41636 13804 41646 13860
rect 44594 13804 44604 13860
rect 44660 13804 45500 13860
rect 45556 13804 45566 13860
rect 51090 13804 51100 13860
rect 51156 13804 55468 13860
rect 55524 13804 55534 13860
rect 5058 13692 5068 13748
rect 5124 13692 6188 13748
rect 6244 13692 6254 13748
rect 7980 13692 16324 13748
rect 17938 13692 17948 13748
rect 18004 13692 21084 13748
rect 21140 13692 21150 13748
rect 25330 13692 25340 13748
rect 25396 13692 26124 13748
rect 26180 13692 26684 13748
rect 26740 13692 26750 13748
rect 27794 13692 27804 13748
rect 27860 13692 42028 13748
rect 42084 13692 42094 13748
rect 45714 13692 45724 13748
rect 45780 13692 47852 13748
rect 47908 13692 49084 13748
rect 49140 13692 50316 13748
rect 50372 13692 50382 13748
rect 54674 13692 54684 13748
rect 54740 13692 54750 13748
rect 55346 13692 55356 13748
rect 55412 13692 55692 13748
rect 55748 13692 55758 13748
rect 1922 13580 1932 13636
rect 1988 13580 2380 13636
rect 2436 13580 2446 13636
rect 8082 13580 8092 13636
rect 8148 13580 9660 13636
rect 9716 13580 9726 13636
rect 10658 13580 10668 13636
rect 10724 13580 12124 13636
rect 12180 13580 12190 13636
rect 14802 13580 14812 13636
rect 14868 13580 15428 13636
rect 24658 13580 24668 13636
rect 24724 13580 26908 13636
rect 26964 13580 26974 13636
rect 27906 13580 27916 13636
rect 27972 13580 28700 13636
rect 28756 13580 29708 13636
rect 29764 13580 29774 13636
rect 34738 13580 34748 13636
rect 34804 13580 35868 13636
rect 35924 13580 37996 13636
rect 38052 13580 38062 13636
rect 38434 13580 38444 13636
rect 38500 13580 40124 13636
rect 40180 13580 41244 13636
rect 41300 13580 41310 13636
rect 15372 13524 15428 13580
rect 3042 13468 3052 13524
rect 3108 13468 3500 13524
rect 3556 13468 3566 13524
rect 8754 13468 8764 13524
rect 8820 13468 15204 13524
rect 15362 13468 15372 13524
rect 15428 13468 15438 13524
rect 16482 13468 16492 13524
rect 16548 13468 22204 13524
rect 22260 13468 23212 13524
rect 23268 13468 23278 13524
rect 24322 13468 24332 13524
rect 24388 13468 26460 13524
rect 26516 13468 26526 13524
rect 34962 13468 34972 13524
rect 35028 13468 35756 13524
rect 35812 13468 37436 13524
rect 37492 13468 37502 13524
rect 39218 13468 39228 13524
rect 39284 13468 39564 13524
rect 39620 13468 39630 13524
rect 41010 13468 41020 13524
rect 41076 13468 42252 13524
rect 42308 13468 42318 13524
rect 48738 13468 48748 13524
rect 48804 13468 49420 13524
rect 49476 13468 49486 13524
rect 51202 13468 51212 13524
rect 51268 13468 53116 13524
rect 53172 13468 53182 13524
rect 15148 13412 15204 13468
rect 54684 13412 54740 13692
rect 2930 13356 2940 13412
rect 2996 13356 3836 13412
rect 3892 13356 3902 13412
rect 6066 13356 6076 13412
rect 6132 13356 6972 13412
rect 7028 13356 7038 13412
rect 10770 13356 10780 13412
rect 10836 13356 11340 13412
rect 11396 13356 11406 13412
rect 15148 13356 21420 13412
rect 21476 13356 21486 13412
rect 54684 13356 58044 13412
rect 58100 13356 58110 13412
rect 8355 13300 8365 13356
rect 8421 13300 8469 13356
rect 8525 13300 8573 13356
rect 8629 13300 8639 13356
rect 22662 13300 22672 13356
rect 22728 13300 22776 13356
rect 22832 13300 22880 13356
rect 22936 13300 22946 13356
rect 36969 13300 36979 13356
rect 37035 13300 37083 13356
rect 37139 13300 37187 13356
rect 37243 13300 37253 13356
rect 51276 13300 51286 13356
rect 51342 13300 51390 13356
rect 51446 13300 51494 13356
rect 51550 13300 51560 13356
rect 14690 13244 14700 13300
rect 14756 13244 15036 13300
rect 15092 13244 15102 13300
rect 29148 13244 33572 13300
rect 29148 13188 29204 13244
rect 33516 13188 33572 13244
rect 1250 13132 1260 13188
rect 1316 13132 22092 13188
rect 22148 13132 22988 13188
rect 23044 13132 23772 13188
rect 23828 13132 25228 13188
rect 25284 13132 27244 13188
rect 27300 13132 27310 13188
rect 28242 13132 28252 13188
rect 28308 13132 28318 13188
rect 29138 13132 29148 13188
rect 29204 13132 29214 13188
rect 30930 13132 30940 13188
rect 30996 13132 33068 13188
rect 33124 13132 33134 13188
rect 33516 13132 46732 13188
rect 46788 13132 47292 13188
rect 47348 13132 47358 13188
rect 48486 13132 48524 13188
rect 48580 13132 48590 13188
rect 50194 13132 50204 13188
rect 50260 13132 51660 13188
rect 51716 13132 52668 13188
rect 52724 13132 54908 13188
rect 54964 13132 55692 13188
rect 55748 13132 56028 13188
rect 56084 13132 56094 13188
rect 57250 13132 57260 13188
rect 57316 13132 57326 13188
rect 28252 13076 28308 13132
rect 57260 13076 57316 13132
rect 59200 13076 60000 13104
rect 1474 13020 1484 13076
rect 1540 13020 5964 13076
rect 6020 13020 6030 13076
rect 10294 13020 10332 13076
rect 10388 13020 10398 13076
rect 11106 13020 11116 13076
rect 11172 13020 12684 13076
rect 12740 13020 12750 13076
rect 17042 13020 17052 13076
rect 17108 13020 19292 13076
rect 19348 13020 19358 13076
rect 19730 13020 19740 13076
rect 19796 13020 20636 13076
rect 20692 13020 22540 13076
rect 22596 13020 23324 13076
rect 23380 13020 23390 13076
rect 28252 13020 45164 13076
rect 45220 13020 45230 13076
rect 51426 13020 51436 13076
rect 51492 13020 53564 13076
rect 53620 13020 53630 13076
rect 53778 13020 53788 13076
rect 53844 13020 55468 13076
rect 55524 13020 55534 13076
rect 55794 13020 55804 13076
rect 55860 13020 56700 13076
rect 56756 13020 56766 13076
rect 57260 13020 60000 13076
rect 59200 12992 60000 13020
rect 4274 12908 4284 12964
rect 4340 12908 4732 12964
rect 4788 12908 4798 12964
rect 16594 12908 16604 12964
rect 16660 12908 17388 12964
rect 17444 12908 18620 12964
rect 18676 12908 18686 12964
rect 20178 12908 20188 12964
rect 20244 12908 21868 12964
rect 21924 12908 21934 12964
rect 30706 12908 30716 12964
rect 30772 12908 31052 12964
rect 31108 12908 31388 12964
rect 31444 12908 31454 12964
rect 37762 12908 37772 12964
rect 37828 12908 40348 12964
rect 40404 12908 40414 12964
rect 44930 12908 44940 12964
rect 44996 12908 45500 12964
rect 45556 12908 45566 12964
rect 48066 12908 48076 12964
rect 48132 12908 48524 12964
rect 48580 12908 48590 12964
rect 50978 12908 50988 12964
rect 51044 12908 51324 12964
rect 51380 12908 52556 12964
rect 52612 12908 53676 12964
rect 53732 12908 54460 12964
rect 54516 12908 54526 12964
rect 55122 12908 55132 12964
rect 55188 12908 56476 12964
rect 56532 12908 56542 12964
rect 1922 12796 1932 12852
rect 1988 12796 2156 12852
rect 2212 12796 2222 12852
rect 9426 12796 9436 12852
rect 9492 12796 15148 12852
rect 18162 12796 18172 12852
rect 18228 12796 18508 12852
rect 18564 12796 18574 12852
rect 30594 12796 30604 12852
rect 30660 12796 32956 12852
rect 33012 12796 33852 12852
rect 33908 12796 33918 12852
rect 35074 12796 35084 12852
rect 35140 12796 35756 12852
rect 35812 12796 35822 12852
rect 38612 12796 51548 12852
rect 51604 12796 51996 12852
rect 52052 12796 52062 12852
rect 53218 12796 53228 12852
rect 53284 12796 57932 12852
rect 57988 12796 57998 12852
rect 15092 12740 15148 12796
rect 38612 12740 38668 12796
rect 3938 12684 3948 12740
rect 4004 12684 7196 12740
rect 7252 12684 7262 12740
rect 15092 12684 19964 12740
rect 20020 12684 20030 12740
rect 34962 12684 34972 12740
rect 35028 12684 35868 12740
rect 35924 12684 35934 12740
rect 36418 12684 36428 12740
rect 36484 12684 38668 12740
rect 41916 12684 45836 12740
rect 45892 12684 45902 12740
rect 47058 12684 47068 12740
rect 47124 12684 47516 12740
rect 47572 12684 47582 12740
rect 53330 12684 53340 12740
rect 53396 12684 54012 12740
rect 54068 12684 54078 12740
rect 55430 12684 55468 12740
rect 55524 12684 55534 12740
rect 56018 12684 56028 12740
rect 56084 12684 57148 12740
rect 57204 12684 57214 12740
rect 41916 12628 41972 12684
rect 32050 12572 32060 12628
rect 32116 12572 41972 12628
rect 55878 12572 55916 12628
rect 55972 12572 55982 12628
rect 15508 12516 15518 12572
rect 15574 12516 15622 12572
rect 15678 12516 15726 12572
rect 15782 12516 15792 12572
rect 29815 12516 29825 12572
rect 29881 12516 29929 12572
rect 29985 12516 30033 12572
rect 30089 12516 30099 12572
rect 44122 12516 44132 12572
rect 44188 12516 44236 12572
rect 44292 12516 44340 12572
rect 44396 12516 44406 12572
rect 58429 12516 58439 12572
rect 58495 12516 58543 12572
rect 58599 12516 58647 12572
rect 58703 12516 58713 12572
rect 3154 12460 3164 12516
rect 3220 12460 3388 12516
rect 37650 12460 37660 12516
rect 37716 12460 38668 12516
rect 38724 12460 38734 12516
rect 48486 12460 48524 12516
rect 48580 12460 48590 12516
rect 3332 12404 3388 12460
rect 3332 12348 6748 12404
rect 6804 12348 6814 12404
rect 9650 12348 9660 12404
rect 9716 12348 10444 12404
rect 10500 12348 11004 12404
rect 11060 12348 11676 12404
rect 11732 12348 12236 12404
rect 12292 12348 13580 12404
rect 13636 12348 13646 12404
rect 14354 12348 14364 12404
rect 14420 12348 16380 12404
rect 16436 12348 16446 12404
rect 18498 12348 18508 12404
rect 18564 12348 18844 12404
rect 18900 12348 18910 12404
rect 23090 12348 23100 12404
rect 23156 12348 23996 12404
rect 24052 12348 24668 12404
rect 24724 12348 25564 12404
rect 25620 12348 26236 12404
rect 26292 12348 26460 12404
rect 26516 12348 27692 12404
rect 27748 12348 28252 12404
rect 28308 12348 28318 12404
rect 34962 12348 34972 12404
rect 35028 12348 35980 12404
rect 36036 12348 36046 12404
rect 42690 12348 42700 12404
rect 42756 12348 44380 12404
rect 44436 12348 45164 12404
rect 45220 12348 45230 12404
rect 47506 12348 47516 12404
rect 47572 12348 47852 12404
rect 47908 12348 49644 12404
rect 49700 12348 50092 12404
rect 50148 12348 50158 12404
rect 54898 12348 54908 12404
rect 54964 12348 55356 12404
rect 55412 12348 55422 12404
rect 56690 12348 56700 12404
rect 56756 12348 57484 12404
rect 57540 12348 58156 12404
rect 58212 12348 58222 12404
rect 4834 12236 4844 12292
rect 4900 12236 18284 12292
rect 18340 12236 18350 12292
rect 32946 12236 32956 12292
rect 33012 12236 35084 12292
rect 35140 12236 35150 12292
rect 47282 12236 47292 12292
rect 47348 12236 48300 12292
rect 48356 12236 48366 12292
rect 49644 12236 51660 12292
rect 51716 12236 52108 12292
rect 52164 12236 52174 12292
rect 55682 12236 55692 12292
rect 55748 12236 57708 12292
rect 57764 12236 57774 12292
rect 0 12180 800 12208
rect 0 12124 2156 12180
rect 2212 12124 2222 12180
rect 3378 12124 3388 12180
rect 3444 12124 3948 12180
rect 4004 12124 4014 12180
rect 8978 12124 8988 12180
rect 9044 12124 10668 12180
rect 10724 12124 10734 12180
rect 19170 12124 19180 12180
rect 19236 12124 19246 12180
rect 21644 12124 23100 12180
rect 23156 12124 23166 12180
rect 28354 12124 28364 12180
rect 28420 12124 29260 12180
rect 29316 12124 29326 12180
rect 33506 12124 33516 12180
rect 33572 12124 34188 12180
rect 34244 12124 35308 12180
rect 35364 12124 35374 12180
rect 48626 12124 48636 12180
rect 48692 12124 49420 12180
rect 49476 12124 49486 12180
rect 0 12096 800 12124
rect 19180 12068 19236 12124
rect 21644 12068 21700 12124
rect 49644 12068 49700 12236
rect 49970 12124 49980 12180
rect 50036 12124 51100 12180
rect 51156 12124 51166 12180
rect 54786 12124 54796 12180
rect 54852 12124 57932 12180
rect 57988 12124 57998 12180
rect 2044 12012 2828 12068
rect 2884 12012 2894 12068
rect 9538 12012 9548 12068
rect 9604 12012 17612 12068
rect 17668 12012 21644 12068
rect 21700 12012 21710 12068
rect 21970 12012 21980 12068
rect 22036 12012 26908 12068
rect 27878 12012 27916 12068
rect 27972 12012 27982 12068
rect 35410 12012 35420 12068
rect 35476 12012 38332 12068
rect 38388 12012 38398 12068
rect 45490 12012 45500 12068
rect 45556 12012 49700 12068
rect 51538 12012 51548 12068
rect 51604 12012 58156 12068
rect 58212 12012 58222 12068
rect 2044 11396 2100 12012
rect 26852 11956 26908 12012
rect 2258 11900 2268 11956
rect 2324 11900 4844 11956
rect 4900 11900 4910 11956
rect 7298 11900 7308 11956
rect 7364 11900 14812 11956
rect 14868 11900 14878 11956
rect 16930 11900 16940 11956
rect 16996 11900 18900 11956
rect 22194 11900 22204 11956
rect 22260 11900 23436 11956
rect 23492 11900 23502 11956
rect 26852 11900 46452 11956
rect 48290 11900 48300 11956
rect 48356 11900 49084 11956
rect 49140 11900 49150 11956
rect 53778 11900 53788 11956
rect 53844 11900 55020 11956
rect 55076 11900 55086 11956
rect 55234 11900 55244 11956
rect 55300 11900 56700 11956
rect 56756 11900 57876 11956
rect 18844 11844 18900 11900
rect 2930 11788 2940 11844
rect 2996 11788 5852 11844
rect 5908 11788 5918 11844
rect 8754 11788 8764 11844
rect 8820 11788 9660 11844
rect 9716 11788 10108 11844
rect 10164 11788 12124 11844
rect 12180 11788 12684 11844
rect 12740 11788 14588 11844
rect 14644 11788 14654 11844
rect 14914 11788 14924 11844
rect 14980 11788 18060 11844
rect 18116 11788 18126 11844
rect 18834 11788 18844 11844
rect 18900 11788 18910 11844
rect 36092 11788 36484 11844
rect 42914 11788 42924 11844
rect 42980 11788 44716 11844
rect 44772 11788 44782 11844
rect 8355 11732 8365 11788
rect 8421 11732 8469 11788
rect 8525 11732 8573 11788
rect 8629 11732 8639 11788
rect 22662 11732 22672 11788
rect 22728 11732 22776 11788
rect 22832 11732 22880 11788
rect 22936 11732 22946 11788
rect 36092 11732 36148 11788
rect 2482 11676 2492 11732
rect 2548 11676 4172 11732
rect 4228 11676 5740 11732
rect 5796 11676 6300 11732
rect 6356 11676 6366 11732
rect 29138 11676 29148 11732
rect 29204 11676 36148 11732
rect 36428 11732 36484 11788
rect 36969 11732 36979 11788
rect 37035 11732 37083 11788
rect 37139 11732 37187 11788
rect 37243 11732 37253 11788
rect 36428 11676 36764 11732
rect 36820 11676 36830 11732
rect 2370 11564 2380 11620
rect 2436 11564 2446 11620
rect 9762 11564 9772 11620
rect 9828 11564 11340 11620
rect 11396 11564 11788 11620
rect 11844 11564 12908 11620
rect 12964 11564 12974 11620
rect 15362 11564 15372 11620
rect 15428 11564 16156 11620
rect 16212 11564 16222 11620
rect 30146 11564 30156 11620
rect 30212 11564 32060 11620
rect 32116 11564 32126 11620
rect 2380 11508 2436 11564
rect 46396 11508 46452 11900
rect 57250 11788 57260 11844
rect 57316 11788 57596 11844
rect 57652 11788 57662 11844
rect 51276 11732 51286 11788
rect 51342 11732 51390 11788
rect 51446 11732 51494 11788
rect 51550 11732 51560 11788
rect 57820 11732 57876 11900
rect 47506 11676 47516 11732
rect 47572 11676 49084 11732
rect 49140 11676 49868 11732
rect 49924 11676 49934 11732
rect 53218 11676 53228 11732
rect 53284 11676 53900 11732
rect 53956 11676 53966 11732
rect 57810 11676 57820 11732
rect 57876 11676 57886 11732
rect 50754 11564 50764 11620
rect 50820 11564 53116 11620
rect 53172 11564 53564 11620
rect 53620 11564 53630 11620
rect 2380 11452 3948 11508
rect 4004 11452 4014 11508
rect 12562 11452 12572 11508
rect 12628 11452 13020 11508
rect 13076 11452 13692 11508
rect 13748 11452 13758 11508
rect 14130 11452 14140 11508
rect 14196 11452 15260 11508
rect 15316 11452 15326 11508
rect 30370 11452 30380 11508
rect 30436 11452 36540 11508
rect 36596 11452 36606 11508
rect 36754 11452 36764 11508
rect 36820 11452 45948 11508
rect 46004 11452 46014 11508
rect 46396 11452 50316 11508
rect 50372 11452 51772 11508
rect 51828 11452 51838 11508
rect 54226 11452 54236 11508
rect 54292 11452 55244 11508
rect 55300 11452 55310 11508
rect 14140 11396 14196 11452
rect 2034 11340 2044 11396
rect 2100 11340 2110 11396
rect 3042 11340 3052 11396
rect 3108 11340 4172 11396
rect 4228 11340 8204 11396
rect 8260 11340 9436 11396
rect 9492 11340 14196 11396
rect 20738 11340 20748 11396
rect 20804 11340 22316 11396
rect 22372 11340 53228 11396
rect 53284 11340 53294 11396
rect 55122 11340 55132 11396
rect 55188 11340 55916 11396
rect 55972 11340 55982 11396
rect 23090 11228 23100 11284
rect 23156 11228 25228 11284
rect 25284 11228 25294 11284
rect 25778 11228 25788 11284
rect 25844 11228 26796 11284
rect 26852 11228 26862 11284
rect 28588 11228 30044 11284
rect 30100 11228 30110 11284
rect 30604 11228 43932 11284
rect 43988 11228 44268 11284
rect 44324 11228 44334 11284
rect 45042 11228 45052 11284
rect 45108 11228 47068 11284
rect 47124 11228 48076 11284
rect 48132 11228 48142 11284
rect 56354 11228 56364 11284
rect 56420 11228 57148 11284
rect 57204 11228 57214 11284
rect 28588 11172 28644 11228
rect 3332 11116 3500 11172
rect 3556 11116 5292 11172
rect 5348 11116 6188 11172
rect 6244 11116 6254 11172
rect 11666 11116 11676 11172
rect 11732 11116 13580 11172
rect 13636 11116 14140 11172
rect 14196 11116 14206 11172
rect 14354 11116 14364 11172
rect 14420 11116 17500 11172
rect 17556 11116 17566 11172
rect 26562 11116 26572 11172
rect 26628 11116 28644 11172
rect 28802 11116 28812 11172
rect 28868 11116 29820 11172
rect 29876 11116 29886 11172
rect 3332 10836 3388 11116
rect 7858 11004 7868 11060
rect 7924 11004 7934 11060
rect 23762 11004 23772 11060
rect 23828 11004 25900 11060
rect 25956 11004 25966 11060
rect 7868 10948 7924 11004
rect 15508 10948 15518 11004
rect 15574 10948 15622 11004
rect 15678 10948 15726 11004
rect 15782 10948 15792 11004
rect 29815 10948 29825 11004
rect 29881 10948 29929 11004
rect 29985 10948 30033 11004
rect 30089 10948 30099 11004
rect 3938 10892 3948 10948
rect 4004 10892 5516 10948
rect 5572 10892 5582 10948
rect 7868 10892 9660 10948
rect 9716 10892 15260 10948
rect 15316 10892 15326 10948
rect 2258 10780 2268 10836
rect 2324 10780 3388 10836
rect 4022 10780 4060 10836
rect 4116 10780 4126 10836
rect 8306 10780 8316 10836
rect 8372 10780 24668 10836
rect 24724 10780 24734 10836
rect 26572 10780 26908 10836
rect 29474 10780 29484 10836
rect 29540 10780 29932 10836
rect 29988 10780 30380 10836
rect 30436 10780 30446 10836
rect 11778 10668 11788 10724
rect 11844 10668 12124 10724
rect 12180 10668 12190 10724
rect 12562 10668 12572 10724
rect 12628 10668 15148 10724
rect 15204 10668 16604 10724
rect 16660 10668 17388 10724
rect 17444 10668 17454 10724
rect 18274 10668 18284 10724
rect 18340 10668 19292 10724
rect 19348 10668 19358 10724
rect 19954 10668 19964 10724
rect 20020 10668 21644 10724
rect 21700 10668 22428 10724
rect 22484 10668 22494 10724
rect 2930 10556 2940 10612
rect 2996 10556 3388 10612
rect 4610 10556 4620 10612
rect 4676 10556 5628 10612
rect 5684 10556 5694 10612
rect 6626 10556 6636 10612
rect 6692 10556 7420 10612
rect 7476 10556 7486 10612
rect 8194 10556 8204 10612
rect 8260 10556 10108 10612
rect 10164 10556 10174 10612
rect 12002 10556 12012 10612
rect 12068 10556 13356 10612
rect 13412 10556 14700 10612
rect 14756 10556 14766 10612
rect 15026 10556 15036 10612
rect 15092 10556 15484 10612
rect 15540 10556 15550 10612
rect 16258 10556 16268 10612
rect 16324 10556 17612 10612
rect 17668 10556 17678 10612
rect 0 10388 800 10416
rect 3332 10388 3388 10556
rect 14700 10500 14756 10556
rect 24668 10500 24724 10780
rect 26572 10612 26628 10780
rect 26852 10724 26908 10780
rect 30604 10724 30660 11228
rect 44268 11172 44324 11228
rect 35186 11116 35196 11172
rect 35252 11116 36316 11172
rect 36372 11116 38220 11172
rect 38276 11116 38286 11172
rect 40226 11116 40236 11172
rect 40292 11116 40684 11172
rect 40740 11116 43596 11172
rect 43652 11116 43662 11172
rect 44268 11116 45276 11172
rect 45332 11116 47964 11172
rect 48020 11116 48030 11172
rect 55458 11116 55468 11172
rect 55524 11116 57372 11172
rect 57428 11116 57438 11172
rect 33170 11004 33180 11060
rect 33236 11004 39900 11060
rect 39956 11004 41692 11060
rect 41748 11004 41758 11060
rect 47012 11004 49644 11060
rect 49700 11004 50652 11060
rect 50708 11004 50718 11060
rect 44122 10948 44132 11004
rect 44188 10948 44236 11004
rect 44292 10948 44340 11004
rect 44396 10948 44406 11004
rect 36530 10892 36540 10948
rect 36596 10892 40404 10948
rect 40348 10836 40404 10892
rect 47012 10836 47068 11004
rect 58429 10948 58439 11004
rect 58495 10948 58543 11004
rect 58599 10948 58647 11004
rect 58703 10948 58713 11004
rect 37762 10780 37772 10836
rect 37828 10780 38332 10836
rect 38388 10780 40124 10836
rect 40180 10780 40190 10836
rect 40348 10780 47068 10836
rect 55458 10780 55468 10836
rect 55524 10780 56252 10836
rect 56308 10780 56318 10836
rect 26852 10668 27132 10724
rect 27188 10668 28476 10724
rect 28532 10668 30660 10724
rect 46386 10668 46396 10724
rect 46452 10668 47852 10724
rect 47908 10668 48860 10724
rect 48916 10668 48926 10724
rect 25442 10556 25452 10612
rect 25508 10556 26572 10612
rect 26628 10556 26638 10612
rect 26786 10556 26796 10612
rect 26852 10556 28812 10612
rect 28868 10556 28878 10612
rect 41906 10556 41916 10612
rect 41972 10556 43036 10612
rect 43092 10556 43102 10612
rect 49634 10556 49644 10612
rect 49700 10556 56924 10612
rect 56980 10556 56990 10612
rect 4946 10444 4956 10500
rect 5012 10444 10556 10500
rect 10612 10444 10622 10500
rect 13020 10444 14364 10500
rect 14420 10444 14430 10500
rect 14700 10444 15372 10500
rect 15428 10444 17052 10500
rect 17108 10444 17118 10500
rect 24668 10444 26908 10500
rect 26964 10444 46284 10500
rect 46340 10444 46620 10500
rect 46676 10444 47068 10500
rect 47124 10444 47404 10500
rect 47460 10444 48636 10500
rect 48692 10444 48702 10500
rect 50418 10444 50428 10500
rect 50484 10444 50652 10500
rect 50708 10444 50718 10500
rect 13020 10388 13076 10444
rect 0 10332 1988 10388
rect 3332 10332 3948 10388
rect 4004 10332 4014 10388
rect 10210 10332 10220 10388
rect 10276 10332 13020 10388
rect 13076 10332 13086 10388
rect 14578 10332 14588 10388
rect 14644 10332 15036 10388
rect 15092 10332 15102 10388
rect 16034 10332 16044 10388
rect 16100 10332 17836 10388
rect 17892 10332 17902 10388
rect 19954 10332 19964 10388
rect 20020 10332 20748 10388
rect 20804 10332 21868 10388
rect 21924 10332 22876 10388
rect 22932 10332 26348 10388
rect 26404 10332 26414 10388
rect 37650 10332 37660 10388
rect 37716 10332 38668 10388
rect 54226 10332 54236 10388
rect 54292 10332 55468 10388
rect 55524 10332 55534 10388
rect 0 10304 800 10332
rect 1932 10276 1988 10332
rect 1922 10220 1932 10276
rect 1988 10220 1998 10276
rect 8355 10164 8365 10220
rect 8421 10164 8469 10220
rect 8525 10164 8573 10220
rect 8629 10164 8639 10220
rect 22662 10164 22672 10220
rect 22728 10164 22776 10220
rect 22832 10164 22880 10220
rect 22936 10164 22946 10220
rect 36969 10164 36979 10220
rect 37035 10164 37083 10220
rect 37139 10164 37187 10220
rect 37243 10164 37253 10220
rect 38612 10164 38668 10332
rect 46956 10220 49308 10276
rect 49364 10220 49374 10276
rect 38612 10108 40348 10164
rect 40404 10108 40414 10164
rect 41020 10108 42420 10164
rect 41020 10052 41076 10108
rect 42364 10052 42420 10108
rect 46956 10052 47012 10220
rect 51276 10164 51286 10220
rect 51342 10164 51390 10220
rect 51446 10164 51494 10220
rect 51550 10164 51560 10220
rect 57922 10108 57932 10164
rect 57988 10108 59332 10164
rect 6066 9996 6076 10052
rect 6132 9996 6860 10052
rect 6916 9996 7756 10052
rect 7812 9996 7822 10052
rect 9090 9996 9100 10052
rect 9156 9996 27356 10052
rect 27412 9996 28364 10052
rect 28420 9996 28430 10052
rect 30706 9996 30716 10052
rect 30772 9996 41076 10052
rect 41234 9996 41244 10052
rect 41300 9996 42140 10052
rect 42196 9996 42206 10052
rect 42364 9996 47012 10052
rect 47954 9996 47964 10052
rect 48020 9996 49980 10052
rect 50036 9996 50046 10052
rect 55234 9996 55244 10052
rect 55300 9996 56700 10052
rect 56756 9996 56766 10052
rect 12786 9884 12796 9940
rect 12852 9884 13692 9940
rect 13748 9884 13758 9940
rect 14242 9884 14252 9940
rect 14308 9884 15148 9940
rect 18274 9884 18284 9940
rect 18340 9884 18956 9940
rect 19012 9884 19022 9940
rect 33730 9884 33740 9940
rect 33796 9884 36428 9940
rect 36484 9884 36494 9940
rect 38434 9884 38444 9940
rect 38500 9884 39788 9940
rect 39844 9884 39854 9940
rect 40114 9884 40124 9940
rect 40180 9884 43372 9940
rect 43428 9884 43438 9940
rect 45154 9884 45164 9940
rect 45220 9884 46956 9940
rect 47012 9884 51660 9940
rect 51716 9884 54684 9940
rect 54740 9884 54750 9940
rect 15092 9828 15148 9884
rect 40124 9828 40180 9884
rect 3042 9772 3052 9828
rect 3108 9772 4508 9828
rect 4564 9772 4574 9828
rect 6290 9772 6300 9828
rect 6356 9772 7084 9828
rect 7140 9772 7150 9828
rect 9090 9772 9100 9828
rect 9156 9772 9884 9828
rect 9940 9772 10444 9828
rect 10500 9772 10510 9828
rect 13794 9772 13804 9828
rect 13860 9772 14476 9828
rect 14532 9772 14542 9828
rect 15092 9772 15708 9828
rect 15764 9772 15774 9828
rect 16146 9772 16156 9828
rect 16212 9772 16828 9828
rect 16884 9772 18060 9828
rect 18116 9772 19180 9828
rect 19236 9772 19246 9828
rect 23314 9772 23324 9828
rect 23380 9772 24444 9828
rect 24500 9772 24510 9828
rect 37762 9772 37772 9828
rect 37828 9772 40180 9828
rect 43474 9772 43484 9828
rect 43540 9772 43550 9828
rect 47618 9772 47628 9828
rect 47684 9772 49532 9828
rect 49588 9772 49598 9828
rect 10444 9716 10500 9772
rect 1922 9660 1932 9716
rect 1988 9660 2604 9716
rect 2660 9660 2670 9716
rect 10444 9660 17836 9716
rect 17892 9660 18844 9716
rect 18900 9660 18910 9716
rect 32834 9660 32844 9716
rect 32900 9660 38108 9716
rect 38164 9660 38174 9716
rect 38322 9660 38332 9716
rect 38388 9660 39340 9716
rect 39396 9660 39406 9716
rect 40898 9660 40908 9716
rect 40964 9660 42364 9716
rect 42420 9660 42430 9716
rect 43484 9604 43540 9772
rect 59276 9716 59332 10108
rect 45266 9660 45276 9716
rect 45332 9660 46508 9716
rect 46564 9660 49868 9716
rect 49924 9660 49934 9716
rect 54898 9660 54908 9716
rect 54964 9660 57372 9716
rect 57428 9660 57438 9716
rect 59052 9660 59332 9716
rect 8082 9548 8092 9604
rect 8148 9548 16268 9604
rect 16324 9548 16334 9604
rect 36418 9548 36428 9604
rect 36484 9548 37100 9604
rect 37156 9548 43540 9604
rect 47618 9548 47628 9604
rect 47684 9548 48412 9604
rect 48468 9548 54572 9604
rect 54628 9548 54638 9604
rect 59052 9492 59108 9660
rect 59200 9492 60000 9520
rect 4498 9436 4508 9492
rect 4564 9436 4844 9492
rect 4900 9436 9828 9492
rect 10098 9436 10108 9492
rect 10164 9436 14812 9492
rect 14868 9436 14878 9492
rect 59052 9436 60000 9492
rect 9772 9380 9828 9436
rect 14812 9380 14868 9436
rect 15508 9380 15518 9436
rect 15574 9380 15622 9436
rect 15678 9380 15726 9436
rect 15782 9380 15792 9436
rect 29815 9380 29825 9436
rect 29881 9380 29929 9436
rect 29985 9380 30033 9436
rect 30089 9380 30099 9436
rect 44122 9380 44132 9436
rect 44188 9380 44236 9436
rect 44292 9380 44340 9436
rect 44396 9380 44406 9436
rect 58429 9380 58439 9436
rect 58495 9380 58543 9436
rect 58599 9380 58647 9436
rect 58703 9380 58713 9436
rect 59200 9408 60000 9436
rect 3602 9324 3612 9380
rect 3668 9324 3836 9380
rect 3892 9324 5068 9380
rect 5124 9324 5134 9380
rect 9762 9324 9772 9380
rect 9828 9324 10668 9380
rect 10724 9324 10734 9380
rect 14690 9324 14700 9380
rect 14756 9324 14868 9380
rect 43474 9324 43484 9380
rect 43540 9324 43550 9380
rect 45378 9324 45388 9380
rect 45444 9324 54348 9380
rect 54404 9324 54414 9380
rect 43484 9268 43540 9324
rect 3378 9212 3388 9268
rect 3444 9212 6300 9268
rect 6356 9212 6366 9268
rect 6738 9212 6748 9268
rect 6804 9212 7532 9268
rect 7588 9212 9660 9268
rect 9716 9212 9726 9268
rect 26852 9212 27468 9268
rect 27524 9212 28028 9268
rect 28084 9212 28094 9268
rect 39442 9212 39452 9268
rect 39508 9212 40012 9268
rect 40068 9212 42812 9268
rect 42868 9212 42878 9268
rect 43484 9212 44716 9268
rect 44772 9212 44782 9268
rect 3836 9156 3892 9212
rect 26852 9156 26908 9212
rect 42588 9156 42644 9212
rect 3826 9100 3836 9156
rect 3892 9100 3902 9156
rect 4498 9100 4508 9156
rect 4564 9100 4844 9156
rect 4900 9100 4910 9156
rect 7746 9100 7756 9156
rect 7812 9100 8988 9156
rect 9044 9100 10668 9156
rect 10724 9100 11228 9156
rect 11284 9100 12572 9156
rect 12628 9100 13804 9156
rect 13860 9100 13870 9156
rect 15586 9100 15596 9156
rect 15652 9100 17724 9156
rect 17780 9100 17790 9156
rect 21074 9100 21084 9156
rect 21140 9100 22540 9156
rect 22596 9100 24556 9156
rect 24612 9100 24622 9156
rect 25778 9100 25788 9156
rect 25844 9100 26684 9156
rect 26740 9100 26908 9156
rect 27346 9100 27356 9156
rect 27412 9100 27422 9156
rect 40450 9100 40460 9156
rect 40516 9100 41580 9156
rect 41636 9100 42028 9156
rect 42084 9100 42094 9156
rect 42578 9100 42588 9156
rect 42644 9100 42654 9156
rect 45266 9100 45276 9156
rect 45332 9100 46732 9156
rect 46788 9100 50428 9156
rect 3490 8988 3500 9044
rect 3556 8988 4060 9044
rect 4116 8988 6076 9044
rect 6132 8988 6142 9044
rect 6514 8988 6524 9044
rect 6580 8988 9996 9044
rect 10052 8988 12012 9044
rect 12068 8988 12078 9044
rect 21970 8988 21980 9044
rect 22036 8988 25452 9044
rect 25508 8988 26124 9044
rect 26180 8988 26190 9044
rect 27356 8932 27412 9100
rect 40908 9044 40964 9100
rect 42028 9044 42084 9100
rect 50372 9044 50428 9100
rect 40898 8988 40908 9044
rect 40964 8988 40974 9044
rect 42028 8988 42812 9044
rect 42868 8988 43036 9044
rect 43092 8988 43102 9044
rect 48178 8988 48188 9044
rect 48244 8988 48972 9044
rect 49028 8988 49038 9044
rect 50372 8988 50764 9044
rect 50820 8988 50830 9044
rect 54786 8988 54796 9044
rect 54852 8988 55356 9044
rect 55412 8988 55422 9044
rect 3378 8876 3388 8932
rect 3444 8876 4956 8932
rect 5012 8876 5022 8932
rect 6626 8876 6636 8932
rect 6692 8876 8540 8932
rect 8596 8876 8606 8932
rect 16706 8876 16716 8932
rect 16772 8876 17836 8932
rect 17892 8876 17902 8932
rect 19618 8876 19628 8932
rect 19684 8876 20412 8932
rect 20468 8876 21308 8932
rect 21364 8876 21374 8932
rect 25666 8876 25676 8932
rect 25732 8876 26572 8932
rect 26628 8876 27412 8932
rect 40226 8876 40236 8932
rect 40292 8876 44604 8932
rect 44660 8876 44670 8932
rect 48738 8876 48748 8932
rect 48804 8876 49980 8932
rect 50036 8876 50046 8932
rect 51314 8876 51324 8932
rect 51380 8876 51772 8932
rect 51828 8876 53564 8932
rect 53620 8876 53630 8932
rect 3938 8764 3948 8820
rect 4004 8764 4396 8820
rect 4452 8764 4462 8820
rect 5170 8764 5180 8820
rect 5236 8764 12908 8820
rect 12964 8764 13356 8820
rect 13412 8764 14476 8820
rect 14532 8764 14924 8820
rect 14980 8764 14990 8820
rect 35186 8764 35196 8820
rect 35252 8764 45500 8820
rect 45556 8764 45566 8820
rect 45938 8764 45948 8820
rect 46004 8764 47516 8820
rect 47572 8764 47582 8820
rect 2482 8652 2492 8708
rect 2548 8652 4844 8708
rect 4900 8652 4910 8708
rect 0 8596 800 8624
rect 8355 8596 8365 8652
rect 8421 8596 8469 8652
rect 8525 8596 8573 8652
rect 8629 8596 8639 8652
rect 22662 8596 22672 8652
rect 22728 8596 22776 8652
rect 22832 8596 22880 8652
rect 22936 8596 22946 8652
rect 36969 8596 36979 8652
rect 37035 8596 37083 8652
rect 37139 8596 37187 8652
rect 37243 8596 37253 8652
rect 51276 8596 51286 8652
rect 51342 8596 51390 8652
rect 51446 8596 51494 8652
rect 51550 8596 51560 8652
rect 0 8540 2716 8596
rect 2772 8540 2782 8596
rect 3826 8540 3836 8596
rect 3892 8540 5404 8596
rect 5460 8540 6860 8596
rect 6916 8540 7644 8596
rect 7700 8540 7710 8596
rect 8866 8540 8876 8596
rect 8932 8540 9660 8596
rect 9716 8540 9726 8596
rect 15474 8540 15484 8596
rect 15540 8540 15932 8596
rect 15988 8540 16380 8596
rect 16436 8540 16446 8596
rect 0 8512 800 8540
rect 4498 8428 4508 8484
rect 4564 8428 18284 8484
rect 18340 8428 18350 8484
rect 26852 8372 26908 8484
rect 26964 8428 26974 8484
rect 31266 8428 31276 8484
rect 31332 8428 33684 8484
rect 37538 8428 37548 8484
rect 37604 8428 40572 8484
rect 40628 8428 40796 8484
rect 40852 8428 40862 8484
rect 54898 8428 54908 8484
rect 54964 8428 56476 8484
rect 56532 8428 56542 8484
rect 33628 8372 33684 8428
rect 3332 8316 3836 8372
rect 3892 8316 3902 8372
rect 4834 8316 4844 8372
rect 4900 8316 5740 8372
rect 5796 8316 5806 8372
rect 10546 8316 10556 8372
rect 10612 8316 26908 8372
rect 28354 8316 28364 8372
rect 28420 8316 31052 8372
rect 31108 8316 31836 8372
rect 31892 8316 33404 8372
rect 33460 8316 33470 8372
rect 33628 8316 36092 8372
rect 36148 8316 36158 8372
rect 41010 8316 41020 8372
rect 41076 8316 41692 8372
rect 41748 8316 42252 8372
rect 42308 8316 42318 8372
rect 52098 8316 52108 8372
rect 52164 8316 53004 8372
rect 53060 8316 54796 8372
rect 54852 8316 54862 8372
rect 3332 8148 3388 8316
rect 3938 8204 3948 8260
rect 4004 8204 6300 8260
rect 6356 8204 6366 8260
rect 7410 8204 7420 8260
rect 7476 8204 8204 8260
rect 8260 8204 8270 8260
rect 9762 8204 9772 8260
rect 9828 8204 10444 8260
rect 10500 8204 10510 8260
rect 11554 8204 11564 8260
rect 11620 8204 12460 8260
rect 12516 8204 13580 8260
rect 13636 8204 15596 8260
rect 15652 8204 15662 8260
rect 20178 8204 20188 8260
rect 20244 8204 21532 8260
rect 21588 8204 21598 8260
rect 21858 8204 21868 8260
rect 21924 8204 23436 8260
rect 23492 8204 23502 8260
rect 24994 8204 25004 8260
rect 25060 8204 25900 8260
rect 25956 8204 25966 8260
rect 26114 8204 26124 8260
rect 26180 8204 26460 8260
rect 26516 8204 26526 8260
rect 27122 8204 27132 8260
rect 27188 8204 29708 8260
rect 29764 8204 29774 8260
rect 31154 8204 31164 8260
rect 31220 8204 32732 8260
rect 32788 8204 32798 8260
rect 38098 8204 38108 8260
rect 38164 8204 39228 8260
rect 39284 8204 39294 8260
rect 41794 8204 41804 8260
rect 41860 8204 42476 8260
rect 42532 8204 43484 8260
rect 43540 8204 43550 8260
rect 45378 8204 45388 8260
rect 45444 8204 45454 8260
rect 48402 8204 48412 8260
rect 48468 8204 48748 8260
rect 48804 8204 48814 8260
rect 52882 8204 52892 8260
rect 52948 8204 55580 8260
rect 55636 8204 55646 8260
rect 2370 8092 2380 8148
rect 2436 8092 3388 8148
rect 3826 8092 3836 8148
rect 3892 8092 6748 8148
rect 6804 8092 6814 8148
rect 7298 8092 7308 8148
rect 7364 8092 7980 8148
rect 8036 8092 8046 8148
rect 8204 8036 8260 8204
rect 45388 8148 45444 8204
rect 9202 8092 9212 8148
rect 9268 8092 10556 8148
rect 10612 8092 11228 8148
rect 11284 8092 11294 8148
rect 14914 8092 14924 8148
rect 14980 8092 15708 8148
rect 15764 8092 15774 8148
rect 20514 8092 20524 8148
rect 20580 8092 25788 8148
rect 25844 8092 25854 8148
rect 26852 8092 29372 8148
rect 29428 8092 29438 8148
rect 32498 8092 32508 8148
rect 32564 8092 33292 8148
rect 33348 8092 33628 8148
rect 33684 8092 33694 8148
rect 34066 8092 34076 8148
rect 34132 8092 34972 8148
rect 35028 8092 35532 8148
rect 35588 8092 35598 8148
rect 38612 8092 45444 8148
rect 26852 8036 26908 8092
rect 38612 8036 38668 8092
rect 2706 7980 2716 8036
rect 2772 7980 4060 8036
rect 4116 7980 4126 8036
rect 8204 7980 10220 8036
rect 10276 7980 10892 8036
rect 10948 7980 10958 8036
rect 25442 7980 25452 8036
rect 25508 7980 26124 8036
rect 26180 7980 26908 8036
rect 33058 7980 33068 8036
rect 33124 7980 34524 8036
rect 34580 7980 35084 8036
rect 35140 7980 35150 8036
rect 35410 7980 35420 8036
rect 35476 7980 38668 8036
rect 45266 7980 45276 8036
rect 45332 7980 46732 8036
rect 46788 7980 46798 8036
rect 48066 7980 48076 8036
rect 48132 7980 55020 8036
rect 55076 7980 55086 8036
rect 5618 7868 5628 7924
rect 5684 7868 13132 7924
rect 13188 7868 13198 7924
rect 23426 7868 23436 7924
rect 23492 7868 25900 7924
rect 25956 7868 26236 7924
rect 26292 7868 26302 7924
rect 15508 7812 15518 7868
rect 15574 7812 15622 7868
rect 15678 7812 15726 7868
rect 15782 7812 15792 7868
rect 29815 7812 29825 7868
rect 29881 7812 29929 7868
rect 29985 7812 30033 7868
rect 30089 7812 30099 7868
rect 44122 7812 44132 7868
rect 44188 7812 44236 7868
rect 44292 7812 44340 7868
rect 44396 7812 44406 7868
rect 58429 7812 58439 7868
rect 58495 7812 58543 7868
rect 58599 7812 58647 7868
rect 58703 7812 58713 7868
rect 2482 7756 2492 7812
rect 2548 7756 3388 7812
rect 3444 7756 7532 7812
rect 7588 7756 7756 7812
rect 7812 7756 7822 7812
rect 2818 7644 2828 7700
rect 2884 7644 8428 7700
rect 8484 7644 8494 7700
rect 12898 7644 12908 7700
rect 12964 7644 13804 7700
rect 13860 7644 13870 7700
rect 24546 7644 24556 7700
rect 24612 7644 27692 7700
rect 27748 7644 27758 7700
rect 12114 7532 12124 7588
rect 12180 7532 13916 7588
rect 13972 7532 13982 7588
rect 25778 7532 25788 7588
rect 25844 7532 30324 7588
rect 34178 7532 34188 7588
rect 34244 7532 35644 7588
rect 35700 7532 35710 7588
rect 41234 7532 41244 7588
rect 41300 7532 42140 7588
rect 42196 7532 42206 7588
rect 43250 7532 43260 7588
rect 43316 7532 45052 7588
rect 45108 7532 45118 7588
rect 57026 7532 57036 7588
rect 57092 7532 57596 7588
rect 57652 7532 57662 7588
rect 30268 7476 30324 7532
rect 2818 7420 2828 7476
rect 2884 7420 3052 7476
rect 3108 7420 3118 7476
rect 4386 7420 4396 7476
rect 4452 7420 6188 7476
rect 6244 7420 6254 7476
rect 11218 7420 11228 7476
rect 11284 7420 11900 7476
rect 11956 7420 14140 7476
rect 14196 7420 14206 7476
rect 18498 7420 18508 7476
rect 18564 7420 19068 7476
rect 19124 7420 20188 7476
rect 20244 7420 20254 7476
rect 21074 7420 21084 7476
rect 21140 7420 28252 7476
rect 28308 7420 28318 7476
rect 28914 7420 28924 7476
rect 28980 7420 29932 7476
rect 29988 7420 29998 7476
rect 30258 7420 30268 7476
rect 30324 7420 30334 7476
rect 32162 7420 32172 7476
rect 32228 7420 34748 7476
rect 34804 7420 34814 7476
rect 40114 7420 40124 7476
rect 40180 7420 41132 7476
rect 41188 7420 42028 7476
rect 42084 7420 42094 7476
rect 44258 7420 44268 7476
rect 44324 7420 46284 7476
rect 46340 7420 46350 7476
rect 57138 7420 57148 7476
rect 57204 7420 58044 7476
rect 58100 7420 58110 7476
rect 28924 7364 28980 7420
rect 27906 7308 27916 7364
rect 27972 7308 28980 7364
rect 33058 7196 33068 7252
rect 33124 7196 33964 7252
rect 34020 7196 34030 7252
rect 2370 7084 2380 7140
rect 2436 7084 3052 7140
rect 3108 7084 3118 7140
rect 14578 7084 14588 7140
rect 14644 7084 15932 7140
rect 15988 7084 15998 7140
rect 8355 7028 8365 7084
rect 8421 7028 8469 7084
rect 8525 7028 8573 7084
rect 8629 7028 8639 7084
rect 22662 7028 22672 7084
rect 22728 7028 22776 7084
rect 22832 7028 22880 7084
rect 22936 7028 22946 7084
rect 36969 7028 36979 7084
rect 37035 7028 37083 7084
rect 37139 7028 37187 7084
rect 37243 7028 37253 7084
rect 51276 7028 51286 7084
rect 51342 7028 51390 7084
rect 51446 7028 51494 7084
rect 51550 7028 51560 7084
rect 31602 6972 31612 7028
rect 31668 6972 31678 7028
rect 31612 6916 31668 6972
rect 23874 6860 23884 6916
rect 23940 6860 24332 6916
rect 24388 6860 25004 6916
rect 25060 6860 30828 6916
rect 30884 6860 31668 6916
rect 43138 6860 43148 6916
rect 43204 6860 43932 6916
rect 43988 6860 44828 6916
rect 44884 6860 44894 6916
rect 52770 6860 52780 6916
rect 52836 6860 57148 6916
rect 57204 6860 57214 6916
rect 0 6804 800 6832
rect 0 6748 1764 6804
rect 4050 6748 4060 6804
rect 4116 6748 4732 6804
rect 4788 6748 4798 6804
rect 16034 6748 16044 6804
rect 16100 6748 17500 6804
rect 17556 6748 18172 6804
rect 18228 6748 18238 6804
rect 18610 6748 18620 6804
rect 18676 6748 20524 6804
rect 20580 6748 21420 6804
rect 21476 6748 21486 6804
rect 26002 6748 26012 6804
rect 26068 6748 30604 6804
rect 30660 6748 30670 6804
rect 39900 6748 43708 6804
rect 43764 6748 43774 6804
rect 45378 6748 45388 6804
rect 45444 6748 53228 6804
rect 53284 6748 53294 6804
rect 0 6720 800 6748
rect 1708 6692 1764 6748
rect 39900 6692 39956 6748
rect 1698 6636 1708 6692
rect 1764 6636 1774 6692
rect 2706 6636 2716 6692
rect 2772 6636 3500 6692
rect 3556 6636 5516 6692
rect 5572 6636 5582 6692
rect 5730 6636 5740 6692
rect 5796 6636 7420 6692
rect 7476 6636 7486 6692
rect 17378 6636 17388 6692
rect 17444 6636 18284 6692
rect 18340 6636 18508 6692
rect 18564 6636 18574 6692
rect 29810 6636 29820 6692
rect 29876 6636 31948 6692
rect 32004 6636 33740 6692
rect 33796 6636 33806 6692
rect 34626 6636 34636 6692
rect 34692 6636 35420 6692
rect 35476 6636 35486 6692
rect 36306 6636 36316 6692
rect 36372 6636 39956 6692
rect 40114 6636 40124 6692
rect 40180 6636 42028 6692
rect 42084 6636 42094 6692
rect 42242 6636 42252 6692
rect 42308 6636 43036 6692
rect 43092 6636 43102 6692
rect 44258 6636 44268 6692
rect 44324 6636 46060 6692
rect 46116 6636 46126 6692
rect 46834 6636 46844 6692
rect 46900 6636 48300 6692
rect 48356 6636 48972 6692
rect 49028 6636 49038 6692
rect 51090 6636 51100 6692
rect 51156 6636 51548 6692
rect 51604 6636 52108 6692
rect 52164 6636 52174 6692
rect 56130 6636 56140 6692
rect 56196 6636 57372 6692
rect 57428 6636 57438 6692
rect 1708 6580 1764 6636
rect 34636 6580 34692 6636
rect 1708 6524 6972 6580
rect 7028 6524 7038 6580
rect 29586 6524 29596 6580
rect 29652 6524 34692 6580
rect 38994 6524 39004 6580
rect 39060 6524 45724 6580
rect 45780 6524 46508 6580
rect 46564 6524 47180 6580
rect 47236 6524 47246 6580
rect 48850 6524 48860 6580
rect 48916 6524 49532 6580
rect 49588 6524 49598 6580
rect 51314 6524 51324 6580
rect 51380 6524 52668 6580
rect 52724 6524 52734 6580
rect 23314 6412 23324 6468
rect 23380 6412 24780 6468
rect 24836 6412 24846 6468
rect 32386 6412 32396 6468
rect 32452 6412 32844 6468
rect 32900 6412 32910 6468
rect 43586 6412 43596 6468
rect 43652 6412 45668 6468
rect 45826 6412 45836 6468
rect 45892 6412 46732 6468
rect 46788 6412 46798 6468
rect 51986 6412 51996 6468
rect 52052 6412 53900 6468
rect 53956 6412 53966 6468
rect 45612 6356 45668 6412
rect 1922 6300 1932 6356
rect 1988 6300 2716 6356
rect 2772 6300 2782 6356
rect 45612 6300 47740 6356
rect 47796 6300 48748 6356
rect 48804 6300 48814 6356
rect 15508 6244 15518 6300
rect 15574 6244 15622 6300
rect 15678 6244 15726 6300
rect 15782 6244 15792 6300
rect 29815 6244 29825 6300
rect 29881 6244 29929 6300
rect 29985 6244 30033 6300
rect 30089 6244 30099 6300
rect 44122 6244 44132 6300
rect 44188 6244 44236 6300
rect 44292 6244 44340 6300
rect 44396 6244 44406 6300
rect 58429 6244 58439 6300
rect 58495 6244 58543 6300
rect 58599 6244 58647 6300
rect 58703 6244 58713 6300
rect 38546 6188 38556 6244
rect 38612 6188 39004 6244
rect 39060 6188 40236 6244
rect 40292 6188 40302 6244
rect 50306 6188 50316 6244
rect 50372 6188 50988 6244
rect 51044 6188 51884 6244
rect 51940 6188 51950 6244
rect 1782 6076 1820 6132
rect 1876 6076 1886 6132
rect 4834 6076 4844 6132
rect 4900 6076 5516 6132
rect 5572 6076 9996 6132
rect 10052 6076 10062 6132
rect 19030 6076 19068 6132
rect 19124 6076 19134 6132
rect 26852 6076 28252 6132
rect 28308 6076 28812 6132
rect 28868 6076 29596 6132
rect 29652 6076 29662 6132
rect 36978 6076 36988 6132
rect 37044 6076 37548 6132
rect 37604 6076 37614 6132
rect 39890 6076 39900 6132
rect 39956 6076 43036 6132
rect 43092 6076 43102 6132
rect 50754 6076 50764 6132
rect 50820 6076 52220 6132
rect 52276 6076 52780 6132
rect 52836 6076 52846 6132
rect 26852 6020 26908 6076
rect 2034 5964 2044 6020
rect 2100 5964 3836 6020
rect 3892 5964 3902 6020
rect 14802 5964 14812 6020
rect 14868 5964 26908 6020
rect 48066 5964 48076 6020
rect 48132 5964 48142 6020
rect 50082 5964 50092 6020
rect 50148 5964 51100 6020
rect 51156 5964 51166 6020
rect 55682 5964 55692 6020
rect 55748 5964 57260 6020
rect 57316 5964 57326 6020
rect 2594 5852 2604 5908
rect 2660 5852 3724 5908
rect 3780 5852 5740 5908
rect 5796 5852 5806 5908
rect 7746 5852 7756 5908
rect 7812 5852 8316 5908
rect 8372 5852 8382 5908
rect 8754 5852 8764 5908
rect 8820 5852 12684 5908
rect 12740 5852 12750 5908
rect 18498 5852 18508 5908
rect 18564 5852 18844 5908
rect 18900 5852 18910 5908
rect 21298 5852 21308 5908
rect 21364 5852 21644 5908
rect 21700 5852 22428 5908
rect 22484 5852 22494 5908
rect 27010 5852 27020 5908
rect 27076 5852 27804 5908
rect 27860 5852 27870 5908
rect 35186 5852 35196 5908
rect 35252 5852 35756 5908
rect 35812 5852 35822 5908
rect 37874 5852 37884 5908
rect 37940 5852 39452 5908
rect 39508 5852 39518 5908
rect 41234 5852 41244 5908
rect 41300 5852 42812 5908
rect 42868 5852 44828 5908
rect 44884 5852 44894 5908
rect 48076 5796 48132 5964
rect 59200 5908 60000 5936
rect 48962 5852 48972 5908
rect 49028 5852 56924 5908
rect 56980 5852 56990 5908
rect 58034 5852 58044 5908
rect 58100 5852 60000 5908
rect 59200 5824 60000 5852
rect 2370 5740 2380 5796
rect 2436 5740 3164 5796
rect 3220 5740 3836 5796
rect 3892 5740 4172 5796
rect 4228 5740 4238 5796
rect 7858 5740 7868 5796
rect 7924 5740 10108 5796
rect 10164 5740 10668 5796
rect 10724 5740 10734 5796
rect 35074 5740 35084 5796
rect 35140 5740 45388 5796
rect 45444 5740 45454 5796
rect 48076 5740 54012 5796
rect 54068 5740 54078 5796
rect 55458 5740 55468 5796
rect 55524 5740 57596 5796
rect 57652 5740 57662 5796
rect 2930 5628 2940 5684
rect 2996 5628 3724 5684
rect 3780 5628 3790 5684
rect 25666 5628 25676 5684
rect 25732 5628 27020 5684
rect 27076 5628 27086 5684
rect 31490 5628 31500 5684
rect 31556 5628 32172 5684
rect 32228 5628 35868 5684
rect 35924 5628 35934 5684
rect 54012 5572 54068 5740
rect 55346 5628 55356 5684
rect 55412 5628 57820 5684
rect 57876 5628 57886 5684
rect 54012 5516 55692 5572
rect 55748 5516 55758 5572
rect 8355 5460 8365 5516
rect 8421 5460 8469 5516
rect 8525 5460 8573 5516
rect 8629 5460 8639 5516
rect 22662 5460 22672 5516
rect 22728 5460 22776 5516
rect 22832 5460 22880 5516
rect 22936 5460 22946 5516
rect 36969 5460 36979 5516
rect 37035 5460 37083 5516
rect 37139 5460 37187 5516
rect 37243 5460 37253 5516
rect 51276 5460 51286 5516
rect 51342 5460 51390 5516
rect 51446 5460 51494 5516
rect 51550 5460 51560 5516
rect 11676 5404 15596 5460
rect 15652 5404 17948 5460
rect 18004 5404 19068 5460
rect 19124 5404 19180 5460
rect 19236 5404 19740 5460
rect 19796 5404 19806 5460
rect 29026 5404 29036 5460
rect 29092 5404 30604 5460
rect 30660 5404 30940 5460
rect 30996 5404 31006 5460
rect 37650 5404 37660 5460
rect 37716 5404 38332 5460
rect 38388 5404 40348 5460
rect 40404 5404 40414 5460
rect 49074 5404 49084 5460
rect 49140 5404 50876 5460
rect 50932 5404 50942 5460
rect 53890 5404 53900 5460
rect 53956 5404 55356 5460
rect 55412 5404 57036 5460
rect 57092 5404 57708 5460
rect 57764 5404 57774 5460
rect 11676 5348 11732 5404
rect 11666 5292 11676 5348
rect 11732 5292 11742 5348
rect 12674 5292 12684 5348
rect 12740 5292 16156 5348
rect 16212 5292 16222 5348
rect 28466 5292 28476 5348
rect 28532 5292 29708 5348
rect 29764 5292 29774 5348
rect 32956 5292 48076 5348
rect 48132 5292 48860 5348
rect 48916 5292 48926 5348
rect 49186 5292 49196 5348
rect 49252 5292 49532 5348
rect 49588 5292 51324 5348
rect 51380 5292 51390 5348
rect 54338 5292 54348 5348
rect 54404 5292 55804 5348
rect 55860 5292 55870 5348
rect 32956 5236 33012 5292
rect 7298 5180 7308 5236
rect 7364 5180 8092 5236
rect 8148 5180 10220 5236
rect 10276 5180 10780 5236
rect 10836 5180 10846 5236
rect 11778 5180 11788 5236
rect 11844 5180 15148 5236
rect 22530 5180 22540 5236
rect 22596 5180 25788 5236
rect 25844 5180 26908 5236
rect 27234 5180 27244 5236
rect 27300 5180 33012 5236
rect 33394 5180 33404 5236
rect 33460 5180 34412 5236
rect 34468 5180 34478 5236
rect 38434 5180 38444 5236
rect 38500 5180 39228 5236
rect 39284 5180 39294 5236
rect 41570 5180 41580 5236
rect 41636 5180 45836 5236
rect 45892 5180 45902 5236
rect 49746 5180 49756 5236
rect 49812 5180 55692 5236
rect 55748 5180 55758 5236
rect 56018 5180 56028 5236
rect 56084 5180 56812 5236
rect 56868 5180 56878 5236
rect 15092 5124 15148 5180
rect 26852 5124 26908 5180
rect 3714 5068 3724 5124
rect 3780 5068 4620 5124
rect 4676 5068 4686 5124
rect 5058 5068 5068 5124
rect 5124 5068 6188 5124
rect 6244 5068 6254 5124
rect 8306 5068 8316 5124
rect 8372 5068 10892 5124
rect 10948 5068 13804 5124
rect 13860 5068 13870 5124
rect 15092 5068 16380 5124
rect 16436 5068 16446 5124
rect 26852 5068 32172 5124
rect 32228 5068 32238 5124
rect 38658 5068 38668 5124
rect 38724 5068 39452 5124
rect 39508 5068 39518 5124
rect 40002 5068 40012 5124
rect 40068 5068 40684 5124
rect 40740 5068 40750 5124
rect 42130 5068 42140 5124
rect 42196 5068 43820 5124
rect 43876 5068 43886 5124
rect 45602 5068 45612 5124
rect 45668 5068 46844 5124
rect 46900 5068 51100 5124
rect 51156 5068 51166 5124
rect 52210 5068 52220 5124
rect 52276 5068 54572 5124
rect 54628 5068 54638 5124
rect 55794 5068 55804 5124
rect 55860 5068 56588 5124
rect 56644 5068 57484 5124
rect 57540 5068 57932 5124
rect 57988 5068 57998 5124
rect 0 5012 800 5040
rect 0 4956 1820 5012
rect 1876 4956 1886 5012
rect 6626 4956 6636 5012
rect 6692 4956 9548 5012
rect 9604 4956 9614 5012
rect 12898 4956 12908 5012
rect 12964 4956 15820 5012
rect 15876 4956 18732 5012
rect 18788 4956 18798 5012
rect 19618 4956 19628 5012
rect 19684 4956 21868 5012
rect 21924 4956 21934 5012
rect 36866 4956 36876 5012
rect 36932 4956 38220 5012
rect 38276 4956 39172 5012
rect 0 4928 800 4956
rect 39116 4900 39172 4956
rect 20626 4844 20636 4900
rect 20692 4844 22876 4900
rect 22932 4844 22942 4900
rect 27122 4844 27132 4900
rect 27188 4844 27468 4900
rect 27524 4844 27534 4900
rect 39106 4844 39116 4900
rect 39172 4844 41916 4900
rect 41972 4844 41982 4900
rect 43932 4844 48972 4900
rect 49028 4844 49644 4900
rect 49700 4844 49710 4900
rect 43932 4788 43988 4844
rect 4162 4732 4172 4788
rect 4228 4732 4956 4788
rect 5012 4732 6076 4788
rect 6132 4732 6142 4788
rect 35410 4732 35420 4788
rect 35476 4732 36092 4788
rect 36148 4732 43988 4788
rect 44930 4732 44940 4788
rect 44996 4732 46732 4788
rect 46788 4732 46798 4788
rect 15508 4676 15518 4732
rect 15574 4676 15622 4732
rect 15678 4676 15726 4732
rect 15782 4676 15792 4732
rect 29815 4676 29825 4732
rect 29881 4676 29929 4732
rect 29985 4676 30033 4732
rect 30089 4676 30099 4732
rect 44122 4676 44132 4732
rect 44188 4676 44236 4732
rect 44292 4676 44340 4732
rect 44396 4676 44406 4732
rect 58429 4676 58439 4732
rect 58495 4676 58543 4732
rect 58599 4676 58647 4732
rect 58703 4676 58713 4732
rect 16706 4620 16716 4676
rect 16772 4620 24556 4676
rect 24612 4620 25228 4676
rect 25284 4620 25294 4676
rect 37426 4620 37436 4676
rect 37492 4620 43708 4676
rect 43764 4620 43774 4676
rect 1810 4508 1820 4564
rect 1876 4508 4396 4564
rect 4452 4508 4462 4564
rect 5170 4508 5180 4564
rect 5236 4508 5628 4564
rect 5684 4508 7196 4564
rect 7252 4508 7262 4564
rect 9762 4508 9772 4564
rect 9828 4508 11004 4564
rect 11060 4508 11070 4564
rect 12786 4508 12796 4564
rect 12852 4508 13468 4564
rect 13524 4508 13534 4564
rect 22082 4508 22092 4564
rect 22148 4508 23996 4564
rect 24052 4508 24062 4564
rect 28690 4508 28700 4564
rect 28756 4508 49868 4564
rect 49924 4508 49934 4564
rect 8194 4396 8204 4452
rect 8260 4396 11788 4452
rect 11844 4396 11854 4452
rect 16370 4396 16380 4452
rect 16436 4396 18060 4452
rect 18116 4396 20076 4452
rect 20132 4396 20142 4452
rect 22754 4396 22764 4452
rect 22820 4396 26684 4452
rect 26740 4396 29372 4452
rect 29428 4396 29438 4452
rect 40338 4396 40348 4452
rect 40404 4396 41356 4452
rect 41412 4396 41422 4452
rect 43922 4396 43932 4452
rect 43988 4396 45164 4452
rect 45220 4396 45230 4452
rect 46722 4396 46732 4452
rect 46788 4396 47404 4452
rect 47460 4396 48860 4452
rect 48916 4396 49308 4452
rect 49364 4396 49374 4452
rect 51538 4396 51548 4452
rect 51604 4396 56924 4452
rect 56980 4396 56990 4452
rect 28588 4340 28644 4396
rect 4722 4284 4732 4340
rect 4788 4284 6300 4340
rect 6356 4284 6366 4340
rect 6850 4284 6860 4340
rect 6916 4284 7532 4340
rect 7588 4284 7598 4340
rect 10658 4284 10668 4340
rect 10724 4284 12012 4340
rect 12068 4284 12078 4340
rect 12450 4284 12460 4340
rect 12516 4284 13356 4340
rect 13412 4284 13422 4340
rect 13906 4284 13916 4340
rect 13972 4284 14476 4340
rect 14532 4284 14542 4340
rect 22418 4284 22428 4340
rect 22484 4284 23772 4340
rect 23828 4284 23838 4340
rect 28578 4284 28588 4340
rect 28644 4284 28654 4340
rect 31154 4284 31164 4340
rect 31220 4284 32284 4340
rect 32340 4284 33068 4340
rect 33124 4284 33134 4340
rect 41570 4284 41580 4340
rect 41636 4284 44156 4340
rect 44212 4284 44222 4340
rect 13916 4228 13972 4284
rect 11442 4172 11452 4228
rect 11508 4172 13132 4228
rect 13188 4172 13972 4228
rect 26460 4172 28364 4228
rect 28420 4172 28924 4228
rect 28980 4172 28990 4228
rect 48066 4172 48076 4228
rect 48132 4172 49532 4228
rect 49588 4172 49598 4228
rect 55906 4172 55916 4228
rect 55972 4172 57932 4228
rect 57988 4172 57998 4228
rect 26460 4116 26516 4172
rect 20962 4060 20972 4116
rect 21028 4060 23436 4116
rect 23492 4060 23502 4116
rect 23762 4060 23772 4116
rect 23828 4060 26460 4116
rect 26516 4060 26526 4116
rect 24098 3948 24108 4004
rect 24164 3948 31948 4004
rect 32004 3948 33292 4004
rect 33348 3948 33358 4004
rect 8355 3892 8365 3948
rect 8421 3892 8469 3948
rect 8525 3892 8573 3948
rect 8629 3892 8639 3948
rect 22662 3892 22672 3948
rect 22728 3892 22776 3948
rect 22832 3892 22880 3948
rect 22936 3892 22946 3948
rect 36969 3892 36979 3948
rect 37035 3892 37083 3948
rect 37139 3892 37187 3948
rect 37243 3892 37253 3948
rect 51276 3892 51286 3948
rect 51342 3892 51390 3948
rect 51446 3892 51494 3948
rect 51550 3892 51560 3948
rect 19058 3724 19068 3780
rect 19124 3724 21868 3780
rect 21924 3724 23660 3780
rect 23716 3724 23726 3780
rect 1810 3612 1820 3668
rect 1876 3612 4732 3668
rect 4788 3612 4798 3668
rect 25666 3612 25676 3668
rect 25732 3612 27356 3668
rect 27412 3612 27422 3668
rect 41346 3612 41356 3668
rect 41412 3612 42364 3668
rect 42420 3612 42430 3668
rect 21074 3500 21084 3556
rect 21140 3500 21644 3556
rect 21700 3500 24668 3556
rect 24724 3500 25452 3556
rect 25508 3500 25518 3556
rect 37538 3500 37548 3556
rect 37604 3500 38108 3556
rect 38164 3500 41132 3556
rect 41188 3500 41468 3556
rect 41524 3500 41534 3556
rect 1698 3388 1708 3444
rect 1764 3388 4284 3444
rect 4340 3388 4350 3444
rect 23762 3388 23772 3444
rect 23828 3388 25788 3444
rect 25844 3388 25854 3444
rect 1810 3276 1820 3332
rect 1876 3276 1886 3332
rect 0 3220 800 3248
rect 1820 3220 1876 3276
rect 0 3164 1876 3220
rect 0 3136 800 3164
rect 15508 3108 15518 3164
rect 15574 3108 15622 3164
rect 15678 3108 15726 3164
rect 15782 3108 15792 3164
rect 29815 3108 29825 3164
rect 29881 3108 29929 3164
rect 29985 3108 30033 3164
rect 30089 3108 30099 3164
rect 44122 3108 44132 3164
rect 44188 3108 44236 3164
rect 44292 3108 44340 3164
rect 44396 3108 44406 3164
rect 58429 3108 58439 3164
rect 58495 3108 58543 3164
rect 58599 3108 58647 3164
rect 58703 3108 58713 3164
rect 56242 2940 56252 2996
rect 56308 2940 59332 2996
rect 59276 2548 59332 2940
rect 59164 2492 59332 2548
rect 59164 2352 59220 2492
rect 59164 2268 60000 2352
rect 59200 2240 60000 2268
rect 0 1428 800 1456
rect 0 1372 1708 1428
rect 1764 1372 1774 1428
rect 0 1344 800 1372
<< via3 >>
rect 15518 26628 15574 26684
rect 15622 26628 15678 26684
rect 15726 26628 15782 26684
rect 29825 26628 29881 26684
rect 29929 26628 29985 26684
rect 30033 26628 30089 26684
rect 44132 26628 44188 26684
rect 44236 26628 44292 26684
rect 44340 26628 44396 26684
rect 58439 26628 58495 26684
rect 58543 26628 58599 26684
rect 58647 26628 58703 26684
rect 26908 26236 26964 26292
rect 8365 25844 8421 25900
rect 8469 25844 8525 25900
rect 8573 25844 8629 25900
rect 22672 25844 22728 25900
rect 22776 25844 22832 25900
rect 22880 25844 22936 25900
rect 36979 25844 37035 25900
rect 37083 25844 37139 25900
rect 37187 25844 37243 25900
rect 51286 25844 51342 25900
rect 51390 25844 51446 25900
rect 51494 25844 51550 25900
rect 15518 25060 15574 25116
rect 15622 25060 15678 25116
rect 15726 25060 15782 25116
rect 29825 25060 29881 25116
rect 29929 25060 29985 25116
rect 30033 25060 30089 25116
rect 44132 25060 44188 25116
rect 44236 25060 44292 25116
rect 44340 25060 44396 25116
rect 58439 25060 58495 25116
rect 58543 25060 58599 25116
rect 58647 25060 58703 25116
rect 8365 24276 8421 24332
rect 8469 24276 8525 24332
rect 8573 24276 8629 24332
rect 22672 24276 22728 24332
rect 22776 24276 22832 24332
rect 22880 24276 22936 24332
rect 36979 24276 37035 24332
rect 37083 24276 37139 24332
rect 37187 24276 37243 24332
rect 51286 24276 51342 24332
rect 51390 24276 51446 24332
rect 51494 24276 51550 24332
rect 15518 23492 15574 23548
rect 15622 23492 15678 23548
rect 15726 23492 15782 23548
rect 29825 23492 29881 23548
rect 29929 23492 29985 23548
rect 30033 23492 30089 23548
rect 44132 23492 44188 23548
rect 44236 23492 44292 23548
rect 44340 23492 44396 23548
rect 58439 23492 58495 23548
rect 58543 23492 58599 23548
rect 58647 23492 58703 23548
rect 16044 22988 16100 23044
rect 26908 22988 26964 23044
rect 8365 22708 8421 22764
rect 8469 22708 8525 22764
rect 8573 22708 8629 22764
rect 22672 22708 22728 22764
rect 22776 22708 22832 22764
rect 22880 22708 22936 22764
rect 36979 22708 37035 22764
rect 37083 22708 37139 22764
rect 37187 22708 37243 22764
rect 51286 22708 51342 22764
rect 51390 22708 51446 22764
rect 51494 22708 51550 22764
rect 16268 22316 16324 22372
rect 15518 21924 15574 21980
rect 15622 21924 15678 21980
rect 15726 21924 15782 21980
rect 29825 21924 29881 21980
rect 29929 21924 29985 21980
rect 30033 21924 30089 21980
rect 44132 21924 44188 21980
rect 44236 21924 44292 21980
rect 44340 21924 44396 21980
rect 58439 21924 58495 21980
rect 58543 21924 58599 21980
rect 58647 21924 58703 21980
rect 16268 21756 16324 21812
rect 8365 21140 8421 21196
rect 8469 21140 8525 21196
rect 8573 21140 8629 21196
rect 22672 21140 22728 21196
rect 22776 21140 22832 21196
rect 22880 21140 22936 21196
rect 36979 21140 37035 21196
rect 37083 21140 37139 21196
rect 37187 21140 37243 21196
rect 51286 21140 51342 21196
rect 51390 21140 51446 21196
rect 51494 21140 51550 21196
rect 1820 21084 1876 21140
rect 16604 20748 16660 20804
rect 15518 20356 15574 20412
rect 15622 20356 15678 20412
rect 15726 20356 15782 20412
rect 29825 20356 29881 20412
rect 29929 20356 29985 20412
rect 30033 20356 30089 20412
rect 44132 20356 44188 20412
rect 44236 20356 44292 20412
rect 44340 20356 44396 20412
rect 58439 20356 58495 20412
rect 58543 20356 58599 20412
rect 58647 20356 58703 20412
rect 38332 20076 38388 20132
rect 38332 19852 38388 19908
rect 8365 19572 8421 19628
rect 8469 19572 8525 19628
rect 8573 19572 8629 19628
rect 22672 19572 22728 19628
rect 22776 19572 22832 19628
rect 22880 19572 22936 19628
rect 36979 19572 37035 19628
rect 37083 19572 37139 19628
rect 37187 19572 37243 19628
rect 51286 19572 51342 19628
rect 51390 19572 51446 19628
rect 51494 19572 51550 19628
rect 15518 18788 15574 18844
rect 15622 18788 15678 18844
rect 15726 18788 15782 18844
rect 29825 18788 29881 18844
rect 29929 18788 29985 18844
rect 30033 18788 30089 18844
rect 44132 18788 44188 18844
rect 44236 18788 44292 18844
rect 44340 18788 44396 18844
rect 58439 18788 58495 18844
rect 58543 18788 58599 18844
rect 58647 18788 58703 18844
rect 27356 18284 27412 18340
rect 8365 18004 8421 18060
rect 8469 18004 8525 18060
rect 8573 18004 8629 18060
rect 22672 18004 22728 18060
rect 22776 18004 22832 18060
rect 22880 18004 22936 18060
rect 36979 18004 37035 18060
rect 37083 18004 37139 18060
rect 37187 18004 37243 18060
rect 27916 17836 27972 17892
rect 51286 18004 51342 18060
rect 51390 18004 51446 18060
rect 51494 18004 51550 18060
rect 15518 17220 15574 17276
rect 15622 17220 15678 17276
rect 15726 17220 15782 17276
rect 29825 17220 29881 17276
rect 29929 17220 29985 17276
rect 30033 17220 30089 17276
rect 44132 17220 44188 17276
rect 44236 17220 44292 17276
rect 44340 17220 44396 17276
rect 58439 17220 58495 17276
rect 58543 17220 58599 17276
rect 58647 17220 58703 17276
rect 8365 16436 8421 16492
rect 8469 16436 8525 16492
rect 8573 16436 8629 16492
rect 22672 16436 22728 16492
rect 22776 16436 22832 16492
rect 22880 16436 22936 16492
rect 36979 16436 37035 16492
rect 37083 16436 37139 16492
rect 37187 16436 37243 16492
rect 51286 16436 51342 16492
rect 51390 16436 51446 16492
rect 51494 16436 51550 16492
rect 27356 16044 27412 16100
rect 50428 15820 50484 15876
rect 15518 15652 15574 15708
rect 15622 15652 15678 15708
rect 15726 15652 15782 15708
rect 29825 15652 29881 15708
rect 29929 15652 29985 15708
rect 30033 15652 30089 15708
rect 44132 15652 44188 15708
rect 44236 15652 44292 15708
rect 44340 15652 44396 15708
rect 58439 15652 58495 15708
rect 58543 15652 58599 15708
rect 58647 15652 58703 15708
rect 50428 15148 50484 15204
rect 8365 14868 8421 14924
rect 8469 14868 8525 14924
rect 8573 14868 8629 14924
rect 22672 14868 22728 14924
rect 22776 14868 22832 14924
rect 22880 14868 22936 14924
rect 36979 14868 37035 14924
rect 37083 14868 37139 14924
rect 37187 14868 37243 14924
rect 51286 14868 51342 14924
rect 51390 14868 51446 14924
rect 51494 14868 51550 14924
rect 10332 14364 10388 14420
rect 15518 14084 15574 14140
rect 15622 14084 15678 14140
rect 15726 14084 15782 14140
rect 16044 13916 16100 13972
rect 14812 13804 14868 13860
rect 29825 14084 29881 14140
rect 29929 14084 29985 14140
rect 30033 14084 30089 14140
rect 44132 14084 44188 14140
rect 44236 14084 44292 14140
rect 44340 14084 44396 14140
rect 58439 14084 58495 14140
rect 58543 14084 58599 14140
rect 58647 14084 58703 14140
rect 55916 13916 55972 13972
rect 16604 13804 16660 13860
rect 55468 13804 55524 13860
rect 14812 13580 14868 13636
rect 8365 13300 8421 13356
rect 8469 13300 8525 13356
rect 8573 13300 8629 13356
rect 22672 13300 22728 13356
rect 22776 13300 22832 13356
rect 22880 13300 22936 13356
rect 36979 13300 37035 13356
rect 37083 13300 37139 13356
rect 37187 13300 37243 13356
rect 51286 13300 51342 13356
rect 51390 13300 51446 13356
rect 51494 13300 51550 13356
rect 48524 13132 48580 13188
rect 10332 13020 10388 13076
rect 55468 12684 55524 12740
rect 55916 12572 55972 12628
rect 15518 12516 15574 12572
rect 15622 12516 15678 12572
rect 15726 12516 15782 12572
rect 29825 12516 29881 12572
rect 29929 12516 29985 12572
rect 30033 12516 30089 12572
rect 44132 12516 44188 12572
rect 44236 12516 44292 12572
rect 44340 12516 44396 12572
rect 58439 12516 58495 12572
rect 58543 12516 58599 12572
rect 58647 12516 58703 12572
rect 48524 12460 48580 12516
rect 27916 12012 27972 12068
rect 8365 11732 8421 11788
rect 8469 11732 8525 11788
rect 8573 11732 8629 11788
rect 22672 11732 22728 11788
rect 22776 11732 22832 11788
rect 22880 11732 22936 11788
rect 36979 11732 37035 11788
rect 37083 11732 37139 11788
rect 37187 11732 37243 11788
rect 51286 11732 51342 11788
rect 51390 11732 51446 11788
rect 51494 11732 51550 11788
rect 36540 11452 36596 11508
rect 15518 10948 15574 11004
rect 15622 10948 15678 11004
rect 15726 10948 15782 11004
rect 29825 10948 29881 11004
rect 29929 10948 29985 11004
rect 30033 10948 30089 11004
rect 4060 10780 4116 10836
rect 44132 10948 44188 11004
rect 44236 10948 44292 11004
rect 44340 10948 44396 11004
rect 36540 10892 36596 10948
rect 58439 10948 58495 11004
rect 58543 10948 58599 11004
rect 58647 10948 58703 11004
rect 8365 10164 8421 10220
rect 8469 10164 8525 10220
rect 8573 10164 8629 10220
rect 22672 10164 22728 10220
rect 22776 10164 22832 10220
rect 22880 10164 22936 10220
rect 36979 10164 37035 10220
rect 37083 10164 37139 10220
rect 37187 10164 37243 10220
rect 51286 10164 51342 10220
rect 51390 10164 51446 10220
rect 51494 10164 51550 10220
rect 14812 9436 14868 9492
rect 15518 9380 15574 9436
rect 15622 9380 15678 9436
rect 15726 9380 15782 9436
rect 29825 9380 29881 9436
rect 29929 9380 29985 9436
rect 30033 9380 30089 9436
rect 44132 9380 44188 9436
rect 44236 9380 44292 9436
rect 44340 9380 44396 9436
rect 58439 9380 58495 9436
rect 58543 9380 58599 9436
rect 58647 9380 58703 9436
rect 8365 8596 8421 8652
rect 8469 8596 8525 8652
rect 8573 8596 8629 8652
rect 22672 8596 22728 8652
rect 22776 8596 22832 8652
rect 22880 8596 22936 8652
rect 36979 8596 37035 8652
rect 37083 8596 37139 8652
rect 37187 8596 37243 8652
rect 51286 8596 51342 8652
rect 51390 8596 51446 8652
rect 51494 8596 51550 8652
rect 15518 7812 15574 7868
rect 15622 7812 15678 7868
rect 15726 7812 15782 7868
rect 29825 7812 29881 7868
rect 29929 7812 29985 7868
rect 30033 7812 30089 7868
rect 44132 7812 44188 7868
rect 44236 7812 44292 7868
rect 44340 7812 44396 7868
rect 58439 7812 58495 7868
rect 58543 7812 58599 7868
rect 58647 7812 58703 7868
rect 8365 7028 8421 7084
rect 8469 7028 8525 7084
rect 8573 7028 8629 7084
rect 22672 7028 22728 7084
rect 22776 7028 22832 7084
rect 22880 7028 22936 7084
rect 36979 7028 37035 7084
rect 37083 7028 37139 7084
rect 37187 7028 37243 7084
rect 51286 7028 51342 7084
rect 51390 7028 51446 7084
rect 51494 7028 51550 7084
rect 4060 6748 4116 6804
rect 15518 6244 15574 6300
rect 15622 6244 15678 6300
rect 15726 6244 15782 6300
rect 29825 6244 29881 6300
rect 29929 6244 29985 6300
rect 30033 6244 30089 6300
rect 44132 6244 44188 6300
rect 44236 6244 44292 6300
rect 44340 6244 44396 6300
rect 58439 6244 58495 6300
rect 58543 6244 58599 6300
rect 58647 6244 58703 6300
rect 1820 6076 1876 6132
rect 19068 6076 19124 6132
rect 8365 5460 8421 5516
rect 8469 5460 8525 5516
rect 8573 5460 8629 5516
rect 22672 5460 22728 5516
rect 22776 5460 22832 5516
rect 22880 5460 22936 5516
rect 36979 5460 37035 5516
rect 37083 5460 37139 5516
rect 37187 5460 37243 5516
rect 51286 5460 51342 5516
rect 51390 5460 51446 5516
rect 51494 5460 51550 5516
rect 19068 5404 19124 5460
rect 15518 4676 15574 4732
rect 15622 4676 15678 4732
rect 15726 4676 15782 4732
rect 29825 4676 29881 4732
rect 29929 4676 29985 4732
rect 30033 4676 30089 4732
rect 44132 4676 44188 4732
rect 44236 4676 44292 4732
rect 44340 4676 44396 4732
rect 58439 4676 58495 4732
rect 58543 4676 58599 4732
rect 58647 4676 58703 4732
rect 8365 3892 8421 3948
rect 8469 3892 8525 3948
rect 8573 3892 8629 3948
rect 22672 3892 22728 3948
rect 22776 3892 22832 3948
rect 22880 3892 22936 3948
rect 36979 3892 37035 3948
rect 37083 3892 37139 3948
rect 37187 3892 37243 3948
rect 51286 3892 51342 3948
rect 51390 3892 51446 3948
rect 51494 3892 51550 3948
rect 15518 3108 15574 3164
rect 15622 3108 15678 3164
rect 15726 3108 15782 3164
rect 29825 3108 29881 3164
rect 29929 3108 29985 3164
rect 30033 3108 30089 3164
rect 44132 3108 44188 3164
rect 44236 3108 44292 3164
rect 44340 3108 44396 3164
rect 58439 3108 58495 3164
rect 58543 3108 58599 3164
rect 58647 3108 58703 3164
<< metal4 >>
rect 8337 25900 8657 26716
rect 8337 25844 8365 25900
rect 8421 25844 8469 25900
rect 8525 25844 8573 25900
rect 8629 25844 8657 25900
rect 8337 24332 8657 25844
rect 8337 24276 8365 24332
rect 8421 24276 8469 24332
rect 8525 24276 8573 24332
rect 8629 24276 8657 24332
rect 8337 22764 8657 24276
rect 8337 22708 8365 22764
rect 8421 22708 8469 22764
rect 8525 22708 8573 22764
rect 8629 22708 8657 22764
rect 8337 21196 8657 22708
rect 1820 21140 1876 21150
rect 1820 6132 1876 21084
rect 8337 21140 8365 21196
rect 8421 21140 8469 21196
rect 8525 21140 8573 21196
rect 8629 21140 8657 21196
rect 8337 19628 8657 21140
rect 8337 19572 8365 19628
rect 8421 19572 8469 19628
rect 8525 19572 8573 19628
rect 8629 19572 8657 19628
rect 8337 18060 8657 19572
rect 8337 18004 8365 18060
rect 8421 18004 8469 18060
rect 8525 18004 8573 18060
rect 8629 18004 8657 18060
rect 8337 16492 8657 18004
rect 8337 16436 8365 16492
rect 8421 16436 8469 16492
rect 8525 16436 8573 16492
rect 8629 16436 8657 16492
rect 8337 14924 8657 16436
rect 8337 14868 8365 14924
rect 8421 14868 8469 14924
rect 8525 14868 8573 14924
rect 8629 14868 8657 14924
rect 8337 13356 8657 14868
rect 15490 26684 15810 26716
rect 15490 26628 15518 26684
rect 15574 26628 15622 26684
rect 15678 26628 15726 26684
rect 15782 26628 15810 26684
rect 15490 25116 15810 26628
rect 15490 25060 15518 25116
rect 15574 25060 15622 25116
rect 15678 25060 15726 25116
rect 15782 25060 15810 25116
rect 15490 23548 15810 25060
rect 15490 23492 15518 23548
rect 15574 23492 15622 23548
rect 15678 23492 15726 23548
rect 15782 23492 15810 23548
rect 15490 21980 15810 23492
rect 22644 25900 22964 26716
rect 29797 26684 30117 26716
rect 29797 26628 29825 26684
rect 29881 26628 29929 26684
rect 29985 26628 30033 26684
rect 30089 26628 30117 26684
rect 22644 25844 22672 25900
rect 22728 25844 22776 25900
rect 22832 25844 22880 25900
rect 22936 25844 22964 25900
rect 22644 24332 22964 25844
rect 22644 24276 22672 24332
rect 22728 24276 22776 24332
rect 22832 24276 22880 24332
rect 22936 24276 22964 24332
rect 15490 21924 15518 21980
rect 15574 21924 15622 21980
rect 15678 21924 15726 21980
rect 15782 21924 15810 21980
rect 15490 20412 15810 21924
rect 15490 20356 15518 20412
rect 15574 20356 15622 20412
rect 15678 20356 15726 20412
rect 15782 20356 15810 20412
rect 15490 18844 15810 20356
rect 15490 18788 15518 18844
rect 15574 18788 15622 18844
rect 15678 18788 15726 18844
rect 15782 18788 15810 18844
rect 15490 17276 15810 18788
rect 15490 17220 15518 17276
rect 15574 17220 15622 17276
rect 15678 17220 15726 17276
rect 15782 17220 15810 17276
rect 15490 15708 15810 17220
rect 15490 15652 15518 15708
rect 15574 15652 15622 15708
rect 15678 15652 15726 15708
rect 15782 15652 15810 15708
rect 8337 13300 8365 13356
rect 8421 13300 8469 13356
rect 8525 13300 8573 13356
rect 8629 13300 8657 13356
rect 8337 11788 8657 13300
rect 10332 14420 10388 14430
rect 10332 13076 10388 14364
rect 15490 14140 15810 15652
rect 15490 14084 15518 14140
rect 15574 14084 15622 14140
rect 15678 14084 15726 14140
rect 15782 14084 15810 14140
rect 10332 13010 10388 13020
rect 14812 13860 14868 13870
rect 14812 13636 14868 13804
rect 8337 11732 8365 11788
rect 8421 11732 8469 11788
rect 8525 11732 8573 11788
rect 8629 11732 8657 11788
rect 4060 10836 4116 10846
rect 4060 6804 4116 10780
rect 4060 6738 4116 6748
rect 8337 10220 8657 11732
rect 8337 10164 8365 10220
rect 8421 10164 8469 10220
rect 8525 10164 8573 10220
rect 8629 10164 8657 10220
rect 8337 8652 8657 10164
rect 14812 9492 14868 13580
rect 14812 9426 14868 9436
rect 15490 12572 15810 14084
rect 16044 23044 16100 23054
rect 16044 13972 16100 22988
rect 22644 22764 22964 24276
rect 26908 26292 26964 26302
rect 26908 23044 26964 26236
rect 26908 22978 26964 22988
rect 29797 25116 30117 26628
rect 29797 25060 29825 25116
rect 29881 25060 29929 25116
rect 29985 25060 30033 25116
rect 30089 25060 30117 25116
rect 29797 23548 30117 25060
rect 29797 23492 29825 23548
rect 29881 23492 29929 23548
rect 29985 23492 30033 23548
rect 30089 23492 30117 23548
rect 22644 22708 22672 22764
rect 22728 22708 22776 22764
rect 22832 22708 22880 22764
rect 22936 22708 22964 22764
rect 16268 22372 16324 22382
rect 16268 21812 16324 22316
rect 16268 21746 16324 21756
rect 22644 21196 22964 22708
rect 22644 21140 22672 21196
rect 22728 21140 22776 21196
rect 22832 21140 22880 21196
rect 22936 21140 22964 21196
rect 16044 13906 16100 13916
rect 16604 20804 16660 20814
rect 16604 13860 16660 20748
rect 16604 13794 16660 13804
rect 22644 19628 22964 21140
rect 22644 19572 22672 19628
rect 22728 19572 22776 19628
rect 22832 19572 22880 19628
rect 22936 19572 22964 19628
rect 22644 18060 22964 19572
rect 29797 21980 30117 23492
rect 29797 21924 29825 21980
rect 29881 21924 29929 21980
rect 29985 21924 30033 21980
rect 30089 21924 30117 21980
rect 29797 20412 30117 21924
rect 29797 20356 29825 20412
rect 29881 20356 29929 20412
rect 29985 20356 30033 20412
rect 30089 20356 30117 20412
rect 29797 18844 30117 20356
rect 29797 18788 29825 18844
rect 29881 18788 29929 18844
rect 29985 18788 30033 18844
rect 30089 18788 30117 18844
rect 22644 18004 22672 18060
rect 22728 18004 22776 18060
rect 22832 18004 22880 18060
rect 22936 18004 22964 18060
rect 22644 16492 22964 18004
rect 22644 16436 22672 16492
rect 22728 16436 22776 16492
rect 22832 16436 22880 16492
rect 22936 16436 22964 16492
rect 22644 14924 22964 16436
rect 27356 18340 27412 18350
rect 27356 16100 27412 18284
rect 27356 16034 27412 16044
rect 27916 17892 27972 17902
rect 22644 14868 22672 14924
rect 22728 14868 22776 14924
rect 22832 14868 22880 14924
rect 22936 14868 22964 14924
rect 15490 12516 15518 12572
rect 15574 12516 15622 12572
rect 15678 12516 15726 12572
rect 15782 12516 15810 12572
rect 15490 11004 15810 12516
rect 15490 10948 15518 11004
rect 15574 10948 15622 11004
rect 15678 10948 15726 11004
rect 15782 10948 15810 11004
rect 15490 9436 15810 10948
rect 8337 8596 8365 8652
rect 8421 8596 8469 8652
rect 8525 8596 8573 8652
rect 8629 8596 8657 8652
rect 8337 7084 8657 8596
rect 8337 7028 8365 7084
rect 8421 7028 8469 7084
rect 8525 7028 8573 7084
rect 8629 7028 8657 7084
rect 1820 6066 1876 6076
rect 8337 5516 8657 7028
rect 8337 5460 8365 5516
rect 8421 5460 8469 5516
rect 8525 5460 8573 5516
rect 8629 5460 8657 5516
rect 8337 3948 8657 5460
rect 8337 3892 8365 3948
rect 8421 3892 8469 3948
rect 8525 3892 8573 3948
rect 8629 3892 8657 3948
rect 8337 3076 8657 3892
rect 15490 9380 15518 9436
rect 15574 9380 15622 9436
rect 15678 9380 15726 9436
rect 15782 9380 15810 9436
rect 15490 7868 15810 9380
rect 15490 7812 15518 7868
rect 15574 7812 15622 7868
rect 15678 7812 15726 7868
rect 15782 7812 15810 7868
rect 15490 6300 15810 7812
rect 15490 6244 15518 6300
rect 15574 6244 15622 6300
rect 15678 6244 15726 6300
rect 15782 6244 15810 6300
rect 15490 4732 15810 6244
rect 22644 13356 22964 14868
rect 22644 13300 22672 13356
rect 22728 13300 22776 13356
rect 22832 13300 22880 13356
rect 22936 13300 22964 13356
rect 22644 11788 22964 13300
rect 27916 12068 27972 17836
rect 27916 12002 27972 12012
rect 29797 17276 30117 18788
rect 29797 17220 29825 17276
rect 29881 17220 29929 17276
rect 29985 17220 30033 17276
rect 30089 17220 30117 17276
rect 29797 15708 30117 17220
rect 29797 15652 29825 15708
rect 29881 15652 29929 15708
rect 29985 15652 30033 15708
rect 30089 15652 30117 15708
rect 29797 14140 30117 15652
rect 29797 14084 29825 14140
rect 29881 14084 29929 14140
rect 29985 14084 30033 14140
rect 30089 14084 30117 14140
rect 29797 12572 30117 14084
rect 29797 12516 29825 12572
rect 29881 12516 29929 12572
rect 29985 12516 30033 12572
rect 30089 12516 30117 12572
rect 22644 11732 22672 11788
rect 22728 11732 22776 11788
rect 22832 11732 22880 11788
rect 22936 11732 22964 11788
rect 22644 10220 22964 11732
rect 22644 10164 22672 10220
rect 22728 10164 22776 10220
rect 22832 10164 22880 10220
rect 22936 10164 22964 10220
rect 22644 8652 22964 10164
rect 22644 8596 22672 8652
rect 22728 8596 22776 8652
rect 22832 8596 22880 8652
rect 22936 8596 22964 8652
rect 22644 7084 22964 8596
rect 22644 7028 22672 7084
rect 22728 7028 22776 7084
rect 22832 7028 22880 7084
rect 22936 7028 22964 7084
rect 19068 6132 19124 6142
rect 19068 5460 19124 6076
rect 19068 5394 19124 5404
rect 22644 5516 22964 7028
rect 22644 5460 22672 5516
rect 22728 5460 22776 5516
rect 22832 5460 22880 5516
rect 22936 5460 22964 5516
rect 15490 4676 15518 4732
rect 15574 4676 15622 4732
rect 15678 4676 15726 4732
rect 15782 4676 15810 4732
rect 15490 3164 15810 4676
rect 15490 3108 15518 3164
rect 15574 3108 15622 3164
rect 15678 3108 15726 3164
rect 15782 3108 15810 3164
rect 15490 3076 15810 3108
rect 22644 3948 22964 5460
rect 22644 3892 22672 3948
rect 22728 3892 22776 3948
rect 22832 3892 22880 3948
rect 22936 3892 22964 3948
rect 22644 3076 22964 3892
rect 29797 11004 30117 12516
rect 36951 25900 37271 26716
rect 36951 25844 36979 25900
rect 37035 25844 37083 25900
rect 37139 25844 37187 25900
rect 37243 25844 37271 25900
rect 36951 24332 37271 25844
rect 36951 24276 36979 24332
rect 37035 24276 37083 24332
rect 37139 24276 37187 24332
rect 37243 24276 37271 24332
rect 36951 22764 37271 24276
rect 36951 22708 36979 22764
rect 37035 22708 37083 22764
rect 37139 22708 37187 22764
rect 37243 22708 37271 22764
rect 36951 21196 37271 22708
rect 36951 21140 36979 21196
rect 37035 21140 37083 21196
rect 37139 21140 37187 21196
rect 37243 21140 37271 21196
rect 36951 19628 37271 21140
rect 44104 26684 44424 26716
rect 44104 26628 44132 26684
rect 44188 26628 44236 26684
rect 44292 26628 44340 26684
rect 44396 26628 44424 26684
rect 44104 25116 44424 26628
rect 44104 25060 44132 25116
rect 44188 25060 44236 25116
rect 44292 25060 44340 25116
rect 44396 25060 44424 25116
rect 44104 23548 44424 25060
rect 44104 23492 44132 23548
rect 44188 23492 44236 23548
rect 44292 23492 44340 23548
rect 44396 23492 44424 23548
rect 44104 21980 44424 23492
rect 44104 21924 44132 21980
rect 44188 21924 44236 21980
rect 44292 21924 44340 21980
rect 44396 21924 44424 21980
rect 44104 20412 44424 21924
rect 44104 20356 44132 20412
rect 44188 20356 44236 20412
rect 44292 20356 44340 20412
rect 44396 20356 44424 20412
rect 38332 20132 38388 20142
rect 38332 19908 38388 20076
rect 38332 19842 38388 19852
rect 36951 19572 36979 19628
rect 37035 19572 37083 19628
rect 37139 19572 37187 19628
rect 37243 19572 37271 19628
rect 36951 18060 37271 19572
rect 36951 18004 36979 18060
rect 37035 18004 37083 18060
rect 37139 18004 37187 18060
rect 37243 18004 37271 18060
rect 36951 16492 37271 18004
rect 36951 16436 36979 16492
rect 37035 16436 37083 16492
rect 37139 16436 37187 16492
rect 37243 16436 37271 16492
rect 36951 14924 37271 16436
rect 36951 14868 36979 14924
rect 37035 14868 37083 14924
rect 37139 14868 37187 14924
rect 37243 14868 37271 14924
rect 36951 13356 37271 14868
rect 36951 13300 36979 13356
rect 37035 13300 37083 13356
rect 37139 13300 37187 13356
rect 37243 13300 37271 13356
rect 36951 11788 37271 13300
rect 36951 11732 36979 11788
rect 37035 11732 37083 11788
rect 37139 11732 37187 11788
rect 37243 11732 37271 11788
rect 29797 10948 29825 11004
rect 29881 10948 29929 11004
rect 29985 10948 30033 11004
rect 30089 10948 30117 11004
rect 29797 9436 30117 10948
rect 36540 11508 36596 11518
rect 36540 10948 36596 11452
rect 36540 10882 36596 10892
rect 29797 9380 29825 9436
rect 29881 9380 29929 9436
rect 29985 9380 30033 9436
rect 30089 9380 30117 9436
rect 29797 7868 30117 9380
rect 29797 7812 29825 7868
rect 29881 7812 29929 7868
rect 29985 7812 30033 7868
rect 30089 7812 30117 7868
rect 29797 6300 30117 7812
rect 29797 6244 29825 6300
rect 29881 6244 29929 6300
rect 29985 6244 30033 6300
rect 30089 6244 30117 6300
rect 29797 4732 30117 6244
rect 29797 4676 29825 4732
rect 29881 4676 29929 4732
rect 29985 4676 30033 4732
rect 30089 4676 30117 4732
rect 29797 3164 30117 4676
rect 29797 3108 29825 3164
rect 29881 3108 29929 3164
rect 29985 3108 30033 3164
rect 30089 3108 30117 3164
rect 29797 3076 30117 3108
rect 36951 10220 37271 11732
rect 36951 10164 36979 10220
rect 37035 10164 37083 10220
rect 37139 10164 37187 10220
rect 37243 10164 37271 10220
rect 36951 8652 37271 10164
rect 36951 8596 36979 8652
rect 37035 8596 37083 8652
rect 37139 8596 37187 8652
rect 37243 8596 37271 8652
rect 36951 7084 37271 8596
rect 36951 7028 36979 7084
rect 37035 7028 37083 7084
rect 37139 7028 37187 7084
rect 37243 7028 37271 7084
rect 36951 5516 37271 7028
rect 36951 5460 36979 5516
rect 37035 5460 37083 5516
rect 37139 5460 37187 5516
rect 37243 5460 37271 5516
rect 36951 3948 37271 5460
rect 36951 3892 36979 3948
rect 37035 3892 37083 3948
rect 37139 3892 37187 3948
rect 37243 3892 37271 3948
rect 36951 3076 37271 3892
rect 44104 18844 44424 20356
rect 44104 18788 44132 18844
rect 44188 18788 44236 18844
rect 44292 18788 44340 18844
rect 44396 18788 44424 18844
rect 44104 17276 44424 18788
rect 44104 17220 44132 17276
rect 44188 17220 44236 17276
rect 44292 17220 44340 17276
rect 44396 17220 44424 17276
rect 44104 15708 44424 17220
rect 51258 25900 51578 26716
rect 51258 25844 51286 25900
rect 51342 25844 51390 25900
rect 51446 25844 51494 25900
rect 51550 25844 51578 25900
rect 51258 24332 51578 25844
rect 51258 24276 51286 24332
rect 51342 24276 51390 24332
rect 51446 24276 51494 24332
rect 51550 24276 51578 24332
rect 51258 22764 51578 24276
rect 51258 22708 51286 22764
rect 51342 22708 51390 22764
rect 51446 22708 51494 22764
rect 51550 22708 51578 22764
rect 51258 21196 51578 22708
rect 51258 21140 51286 21196
rect 51342 21140 51390 21196
rect 51446 21140 51494 21196
rect 51550 21140 51578 21196
rect 51258 19628 51578 21140
rect 51258 19572 51286 19628
rect 51342 19572 51390 19628
rect 51446 19572 51494 19628
rect 51550 19572 51578 19628
rect 51258 18060 51578 19572
rect 51258 18004 51286 18060
rect 51342 18004 51390 18060
rect 51446 18004 51494 18060
rect 51550 18004 51578 18060
rect 51258 16492 51578 18004
rect 51258 16436 51286 16492
rect 51342 16436 51390 16492
rect 51446 16436 51494 16492
rect 51550 16436 51578 16492
rect 44104 15652 44132 15708
rect 44188 15652 44236 15708
rect 44292 15652 44340 15708
rect 44396 15652 44424 15708
rect 44104 14140 44424 15652
rect 50428 15876 50484 15886
rect 50428 15204 50484 15820
rect 50428 15138 50484 15148
rect 44104 14084 44132 14140
rect 44188 14084 44236 14140
rect 44292 14084 44340 14140
rect 44396 14084 44424 14140
rect 44104 12572 44424 14084
rect 51258 14924 51578 16436
rect 51258 14868 51286 14924
rect 51342 14868 51390 14924
rect 51446 14868 51494 14924
rect 51550 14868 51578 14924
rect 51258 13356 51578 14868
rect 58411 26684 58731 26716
rect 58411 26628 58439 26684
rect 58495 26628 58543 26684
rect 58599 26628 58647 26684
rect 58703 26628 58731 26684
rect 58411 25116 58731 26628
rect 58411 25060 58439 25116
rect 58495 25060 58543 25116
rect 58599 25060 58647 25116
rect 58703 25060 58731 25116
rect 58411 23548 58731 25060
rect 58411 23492 58439 23548
rect 58495 23492 58543 23548
rect 58599 23492 58647 23548
rect 58703 23492 58731 23548
rect 58411 21980 58731 23492
rect 58411 21924 58439 21980
rect 58495 21924 58543 21980
rect 58599 21924 58647 21980
rect 58703 21924 58731 21980
rect 58411 20412 58731 21924
rect 58411 20356 58439 20412
rect 58495 20356 58543 20412
rect 58599 20356 58647 20412
rect 58703 20356 58731 20412
rect 58411 18844 58731 20356
rect 58411 18788 58439 18844
rect 58495 18788 58543 18844
rect 58599 18788 58647 18844
rect 58703 18788 58731 18844
rect 58411 17276 58731 18788
rect 58411 17220 58439 17276
rect 58495 17220 58543 17276
rect 58599 17220 58647 17276
rect 58703 17220 58731 17276
rect 58411 15708 58731 17220
rect 58411 15652 58439 15708
rect 58495 15652 58543 15708
rect 58599 15652 58647 15708
rect 58703 15652 58731 15708
rect 58411 14140 58731 15652
rect 58411 14084 58439 14140
rect 58495 14084 58543 14140
rect 58599 14084 58647 14140
rect 58703 14084 58731 14140
rect 55916 13972 55972 13982
rect 51258 13300 51286 13356
rect 51342 13300 51390 13356
rect 51446 13300 51494 13356
rect 51550 13300 51578 13356
rect 44104 12516 44132 12572
rect 44188 12516 44236 12572
rect 44292 12516 44340 12572
rect 44396 12516 44424 12572
rect 44104 11004 44424 12516
rect 48524 13188 48580 13198
rect 48524 12516 48580 13132
rect 48524 12450 48580 12460
rect 44104 10948 44132 11004
rect 44188 10948 44236 11004
rect 44292 10948 44340 11004
rect 44396 10948 44424 11004
rect 44104 9436 44424 10948
rect 44104 9380 44132 9436
rect 44188 9380 44236 9436
rect 44292 9380 44340 9436
rect 44396 9380 44424 9436
rect 44104 7868 44424 9380
rect 44104 7812 44132 7868
rect 44188 7812 44236 7868
rect 44292 7812 44340 7868
rect 44396 7812 44424 7868
rect 44104 6300 44424 7812
rect 44104 6244 44132 6300
rect 44188 6244 44236 6300
rect 44292 6244 44340 6300
rect 44396 6244 44424 6300
rect 44104 4732 44424 6244
rect 44104 4676 44132 4732
rect 44188 4676 44236 4732
rect 44292 4676 44340 4732
rect 44396 4676 44424 4732
rect 44104 3164 44424 4676
rect 44104 3108 44132 3164
rect 44188 3108 44236 3164
rect 44292 3108 44340 3164
rect 44396 3108 44424 3164
rect 44104 3076 44424 3108
rect 51258 11788 51578 13300
rect 55468 13860 55524 13870
rect 55468 12740 55524 13804
rect 55468 12674 55524 12684
rect 55916 12628 55972 13916
rect 55916 12562 55972 12572
rect 58411 12572 58731 14084
rect 51258 11732 51286 11788
rect 51342 11732 51390 11788
rect 51446 11732 51494 11788
rect 51550 11732 51578 11788
rect 51258 10220 51578 11732
rect 51258 10164 51286 10220
rect 51342 10164 51390 10220
rect 51446 10164 51494 10220
rect 51550 10164 51578 10220
rect 51258 8652 51578 10164
rect 51258 8596 51286 8652
rect 51342 8596 51390 8652
rect 51446 8596 51494 8652
rect 51550 8596 51578 8652
rect 51258 7084 51578 8596
rect 51258 7028 51286 7084
rect 51342 7028 51390 7084
rect 51446 7028 51494 7084
rect 51550 7028 51578 7084
rect 51258 5516 51578 7028
rect 51258 5460 51286 5516
rect 51342 5460 51390 5516
rect 51446 5460 51494 5516
rect 51550 5460 51578 5516
rect 51258 3948 51578 5460
rect 51258 3892 51286 3948
rect 51342 3892 51390 3948
rect 51446 3892 51494 3948
rect 51550 3892 51578 3948
rect 51258 3076 51578 3892
rect 58411 12516 58439 12572
rect 58495 12516 58543 12572
rect 58599 12516 58647 12572
rect 58703 12516 58731 12572
rect 58411 11004 58731 12516
rect 58411 10948 58439 11004
rect 58495 10948 58543 11004
rect 58599 10948 58647 11004
rect 58703 10948 58731 11004
rect 58411 9436 58731 10948
rect 58411 9380 58439 9436
rect 58495 9380 58543 9436
rect 58599 9380 58647 9436
rect 58703 9380 58731 9436
rect 58411 7868 58731 9380
rect 58411 7812 58439 7868
rect 58495 7812 58543 7868
rect 58599 7812 58647 7868
rect 58703 7812 58731 7868
rect 58411 6300 58731 7812
rect 58411 6244 58439 6300
rect 58495 6244 58543 6300
rect 58599 6244 58647 6300
rect 58703 6244 58731 6300
rect 58411 4732 58731 6244
rect 58411 4676 58439 4732
rect 58495 4676 58543 4732
rect 58599 4676 58647 4732
rect 58703 4676 58731 4732
rect 58411 3164 58731 4676
rect 58411 3108 58439 3164
rect 58495 3108 58543 3164
rect 58599 3108 58647 3164
rect 58703 3108 58731 3164
rect 58411 3076 58731 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _0692_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0693_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7392 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _0694_
timestamp 1698431365
transform -1 0 6944 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0695_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 1 25088
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0696_
timestamp 1698431365
transform -1 0 10528 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0697_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0698_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0699_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2352 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0700_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5264 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0701_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5040 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _0702_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2352 0 1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0703_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _0704_
timestamp 1698431365
transform -1 0 8064 0 1 21952
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0705_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__and3_4  _0706_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0707_
timestamp 1698431365
transform 1 0 6944 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0708_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16016 0 1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0709_
timestamp 1698431365
transform -1 0 20384 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0710_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0711_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0712_
timestamp 1698431365
transform 1 0 1904 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _0713_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2800 0 -1 20384
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0714_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0715_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6384 0 1 20384
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0716_
timestamp 1698431365
transform -1 0 12208 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0717_
timestamp 1698431365
transform 1 0 3136 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0718_
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _0719_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6496 0 -1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0720_
timestamp 1698431365
transform -1 0 17472 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0721_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6160 0 -1 14112
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0722_
timestamp 1698431365
transform 1 0 2800 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  _0723_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0724_
timestamp 1698431365
transform -1 0 16800 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0725_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23072 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0726_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0727_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1904 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0728_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4032 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0729_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3024 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0730_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2800 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0731_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9296 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0732_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16016 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _0733_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0734_
timestamp 1698431365
transform 1 0 5488 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0735_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16800 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0736_
timestamp 1698431365
transform 1 0 10976 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0737_
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0738_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0739_
timestamp 1698431365
transform -1 0 8960 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0740_
timestamp 1698431365
transform -1 0 10080 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0741_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0742_
timestamp 1698431365
transform 1 0 13888 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0743_
timestamp 1698431365
transform 1 0 1904 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0744_
timestamp 1698431365
transform 1 0 2688 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0745_
timestamp 1698431365
transform 1 0 8736 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0746_
timestamp 1698431365
transform -1 0 19376 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0747_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0748_
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0749_
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0750_
timestamp 1698431365
transform -1 0 19824 0 -1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0751_
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0752_
timestamp 1698431365
transform -1 0 7392 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0753_
timestamp 1698431365
transform 1 0 6720 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0754_
timestamp 1698431365
transform -1 0 11088 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _0755_
timestamp 1698431365
transform 1 0 8736 0 1 21952
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0756_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0757_
timestamp 1698431365
transform 1 0 6384 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_4  _0758_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 -1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0759_
timestamp 1698431365
transform 1 0 8512 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0760_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0761_
timestamp 1698431365
transform 1 0 6272 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0762_
timestamp 1698431365
transform 1 0 7392 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0763_
timestamp 1698431365
transform 1 0 3472 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0764_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0765_
timestamp 1698431365
transform -1 0 16912 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0766_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12096 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0767_
timestamp 1698431365
transform 1 0 11648 0 -1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0768_
timestamp 1698431365
transform 1 0 10416 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _0769_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0770_
timestamp 1698431365
transform -1 0 13664 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0771_
timestamp 1698431365
transform 1 0 11088 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0772_
timestamp 1698431365
transform -1 0 2800 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0773_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0774_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11872 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0775_
timestamp 1698431365
transform -1 0 15904 0 -1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0776_
timestamp 1698431365
transform -1 0 16352 0 1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0777_
timestamp 1698431365
transform 1 0 11424 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0778_
timestamp 1698431365
transform 1 0 11312 0 -1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0779_
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0780_
timestamp 1698431365
transform -1 0 9520 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0781_
timestamp 1698431365
transform -1 0 15456 0 -1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0782_
timestamp 1698431365
transform 1 0 9520 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0783_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0784_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11424 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0785_
timestamp 1698431365
transform -1 0 11424 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0786_
timestamp 1698431365
transform -1 0 7280 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0787_
timestamp 1698431365
transform -1 0 13328 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0788_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _0789_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0790_
timestamp 1698431365
transform -1 0 9184 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0791_
timestamp 1698431365
transform -1 0 17024 0 -1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0792_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15680 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0793_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0794_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0795_
timestamp 1698431365
transform -1 0 11984 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0796_
timestamp 1698431365
transform 1 0 13888 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0797_
timestamp 1698431365
transform -1 0 22848 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0798_
timestamp 1698431365
transform -1 0 21616 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0799_
timestamp 1698431365
transform 1 0 22624 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0800_
timestamp 1698431365
transform 1 0 20384 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0801_
timestamp 1698431365
transform -1 0 22288 0 -1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0802_
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _0803_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0804_
timestamp 1698431365
transform 1 0 21728 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0805_
timestamp 1698431365
transform 1 0 26320 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0806_
timestamp 1698431365
transform 1 0 26992 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0807_
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _0808_
timestamp 1698431365
transform 1 0 23520 0 1 10976
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0809_
timestamp 1698431365
transform -1 0 31024 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0810_
timestamp 1698431365
transform -1 0 35840 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0811_
timestamp 1698431365
transform -1 0 16016 0 1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0812_
timestamp 1698431365
transform 1 0 12096 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0813_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _0814_
timestamp 1698431365
transform 1 0 15904 0 1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0815_
timestamp 1698431365
transform 1 0 8288 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0816_
timestamp 1698431365
transform -1 0 10976 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0817_
timestamp 1698431365
transform -1 0 16464 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0818_
timestamp 1698431365
transform -1 0 18256 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0819_
timestamp 1698431365
transform 1 0 18256 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0820_
timestamp 1698431365
transform -1 0 21840 0 -1 14112
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0821_
timestamp 1698431365
transform -1 0 19040 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0822_
timestamp 1698431365
transform 1 0 8512 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0823_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0824_
timestamp 1698431365
transform 1 0 13664 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0825_
timestamp 1698431365
transform -1 0 16912 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _0826_
timestamp 1698431365
transform -1 0 19936 0 1 17248
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0827_
timestamp 1698431365
transform -1 0 23072 0 -1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0828_
timestamp 1698431365
transform -1 0 16576 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0829_
timestamp 1698431365
transform 1 0 21840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _0830_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0831_
timestamp 1698431365
transform -1 0 19936 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0832_
timestamp 1698431365
transform -1 0 23632 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0833_
timestamp 1698431365
transform -1 0 22960 0 -1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0834_
timestamp 1698431365
transform -1 0 10192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0835_
timestamp 1698431365
transform 1 0 7392 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0836_
timestamp 1698431365
transform 1 0 16464 0 1 14112
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0837_
timestamp 1698431365
transform 1 0 16800 0 1 15680
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0838_
timestamp 1698431365
transform 1 0 17360 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0839_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0840_
timestamp 1698431365
transform -1 0 16912 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0841_
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _0842_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21952 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0843_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0844_
timestamp 1698431365
transform -1 0 23408 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0845_
timestamp 1698431365
transform -1 0 22848 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0846_
timestamp 1698431365
transform -1 0 26208 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0847_
timestamp 1698431365
transform -1 0 27104 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0848_
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0849_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _0850_
timestamp 1698431365
transform 1 0 23184 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0851_
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0852_
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0853_
timestamp 1698431365
transform -1 0 37408 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _0854_
timestamp 1698431365
transform 1 0 37408 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _0855_
timestamp 1698431365
transform 1 0 21952 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0856_
timestamp 1698431365
transform 1 0 28224 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0857_
timestamp 1698431365
transform -1 0 23184 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0858_
timestamp 1698431365
transform -1 0 30352 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0859_
timestamp 1698431365
transform 1 0 27888 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0860_
timestamp 1698431365
transform -1 0 35392 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0861_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _0862_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0863_
timestamp 1698431365
transform -1 0 29344 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0864_
timestamp 1698431365
transform 1 0 35728 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0865_
timestamp 1698431365
transform 1 0 35952 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0866_
timestamp 1698431365
transform 1 0 37520 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0867_
timestamp 1698431365
transform -1 0 27888 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0868_
timestamp 1698431365
transform -1 0 26880 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0869_
timestamp 1698431365
transform 1 0 26432 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0870_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0871_
timestamp 1698431365
transform 1 0 34272 0 -1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0872_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 -1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0873_
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0874_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0875_
timestamp 1698431365
transform 1 0 34720 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0876_
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0877_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0878_
timestamp 1698431365
transform -1 0 35392 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0879_
timestamp 1698431365
transform -1 0 35280 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0880_
timestamp 1698431365
transform 1 0 34832 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0881_
timestamp 1698431365
transform -1 0 35168 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0882_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0883_
timestamp 1698431365
transform 1 0 31920 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0884_
timestamp 1698431365
transform -1 0 32256 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0885_
timestamp 1698431365
transform 1 0 29008 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _0886_
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0887_
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0888_
timestamp 1698431365
transform 1 0 31024 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0889_
timestamp 1698431365
transform -1 0 31584 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0890_
timestamp 1698431365
transform -1 0 27440 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0891_
timestamp 1698431365
transform -1 0 28784 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0892_
timestamp 1698431365
transform 1 0 24304 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0893_
timestamp 1698431365
transform 1 0 26656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0894_
timestamp 1698431365
transform -1 0 25648 0 1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0895_
timestamp 1698431365
transform 1 0 23520 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0896_
timestamp 1698431365
transform -1 0 26656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0897_
timestamp 1698431365
transform 1 0 27552 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0898_
timestamp 1698431365
transform 1 0 26432 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0899_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27552 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0900_
timestamp 1698431365
transform -1 0 34832 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0901_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26992 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _0902_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30688 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0903_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0904_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0905_
timestamp 1698431365
transform 1 0 35168 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0906_
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0907_
timestamp 1698431365
transform 1 0 25872 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0908_
timestamp 1698431365
transform 1 0 29568 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0909_
timestamp 1698431365
transform -1 0 33376 0 1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0910_
timestamp 1698431365
transform -1 0 34048 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0911_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0912_
timestamp 1698431365
transform -1 0 33936 0 1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0913_
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0914_
timestamp 1698431365
transform -1 0 31920 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _0915_
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0916_
timestamp 1698431365
transform 1 0 31136 0 1 12544
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0917_
timestamp 1698431365
transform 1 0 34048 0 -1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0918_
timestamp 1698431365
transform -1 0 39088 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _0919_
timestamp 1698431365
transform -1 0 42000 0 1 12544
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _0920_
timestamp 1698431365
transform 1 0 36624 0 -1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0921_
timestamp 1698431365
transform -1 0 39536 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0922_
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0923_
timestamp 1698431365
transform 1 0 30240 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0924_
timestamp 1698431365
transform -1 0 35952 0 -1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0925_
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0926_
timestamp 1698431365
transform -1 0 30800 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0927_
timestamp 1698431365
transform 1 0 30016 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _0928_
timestamp 1698431365
transform 1 0 42448 0 1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0929_
timestamp 1698431365
transform 1 0 23072 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0930_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0931_
timestamp 1698431365
transform -1 0 26432 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0932_
timestamp 1698431365
transform -1 0 25760 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0933_
timestamp 1698431365
transform -1 0 22624 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0934_
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0935_
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0936_
timestamp 1698431365
transform -1 0 25872 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0937_
timestamp 1698431365
transform -1 0 26656 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0938_
timestamp 1698431365
transform 1 0 19824 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0939_
timestamp 1698431365
transform 1 0 19824 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0940_
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0941_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0942_
timestamp 1698431365
transform -1 0 24976 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0943_
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0944_
timestamp 1698431365
transform -1 0 24640 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0945_
timestamp 1698431365
transform 1 0 38528 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0946_
timestamp 1698431365
transform 1 0 39536 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0947_
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0948_
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0949_
timestamp 1698431365
transform -1 0 31136 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0950_
timestamp 1698431365
transform 1 0 30912 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0951_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0952_
timestamp 1698431365
transform 1 0 39760 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0953_
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_4  _0954_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34160 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _0955_
timestamp 1698431365
transform -1 0 43232 0 -1 20384
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0956_
timestamp 1698431365
transform 1 0 39984 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0957_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0958_
timestamp 1698431365
transform 1 0 40992 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _0959_
timestamp 1698431365
transform 1 0 41328 0 1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0960_
timestamp 1698431365
transform 1 0 42896 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _0961_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33376 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _0962_
timestamp 1698431365
transform 1 0 41328 0 -1 12544
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0963_
timestamp 1698431365
transform 1 0 42896 0 -1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0964_
timestamp 1698431365
transform -1 0 47600 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0965_
timestamp 1698431365
transform -1 0 41776 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0966_
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0967_
timestamp 1698431365
transform 1 0 27552 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0968_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41776 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0969_
timestamp 1698431365
transform -1 0 6384 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _0970_
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0971_
timestamp 1698431365
transform 1 0 2128 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _0972_
timestamp 1698431365
transform 1 0 2352 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0973_
timestamp 1698431365
transform 1 0 26992 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0974_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0975_
timestamp 1698431365
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0976_
timestamp 1698431365
transform 1 0 48944 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0977_
timestamp 1698431365
transform -1 0 7168 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0978_
timestamp 1698431365
transform -1 0 4928 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _0979_
timestamp 1698431365
transform 1 0 5264 0 -1 10976
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0980_
timestamp 1698431365
transform -1 0 29232 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0981_
timestamp 1698431365
transform 1 0 46256 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0982_
timestamp 1698431365
transform 1 0 46704 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0983_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0984_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44576 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0985_
timestamp 1698431365
transform -1 0 20272 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0986_
timestamp 1698431365
transform 1 0 26208 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0987_
timestamp 1698431365
transform -1 0 51520 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0988_
timestamp 1698431365
transform 1 0 48496 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0989_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30464 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0990_
timestamp 1698431365
transform -1 0 36624 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _0991_
timestamp 1698431365
transform 1 0 37408 0 -1 23520
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0992_
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0993_
timestamp 1698431365
transform -1 0 33600 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0994_
timestamp 1698431365
transform -1 0 35168 0 -1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0995_
timestamp 1698431365
transform 1 0 35616 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0996_
timestamp 1698431365
transform -1 0 36848 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0997_
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0998_
timestamp 1698431365
transform -1 0 39984 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0999_
timestamp 1698431365
transform 1 0 32592 0 1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1000_
timestamp 1698431365
transform 1 0 35840 0 -1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1001_
timestamp 1698431365
transform 1 0 31360 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1002_
timestamp 1698431365
transform -1 0 35728 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1003_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1004_
timestamp 1698431365
transform -1 0 39424 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1005_
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1006_
timestamp 1698431365
transform 1 0 37408 0 1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1007_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42672 0 1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1008_
timestamp 1698431365
transform 1 0 34048 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1009_
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1010_
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1011_
timestamp 1698431365
transform -1 0 29008 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1012_
timestamp 1698431365
transform -1 0 28672 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1013_
timestamp 1698431365
transform -1 0 37408 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  _1014_
timestamp 1698431365
transform 1 0 38080 0 -1 21952
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _1015_
timestamp 1698431365
transform 1 0 42448 0 1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1016_
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1017_
timestamp 1698431365
transform 1 0 22512 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1018_
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1019_
timestamp 1698431365
transform 1 0 22960 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1020_
timestamp 1698431365
transform 1 0 39536 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1021_
timestamp 1698431365
transform -1 0 36624 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1022_
timestamp 1698431365
transform 1 0 41440 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1023_
timestamp 1698431365
transform -1 0 36288 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1024_
timestamp 1698431365
transform 1 0 34944 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1025_
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1026_
timestamp 1698431365
transform -1 0 43904 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1027_
timestamp 1698431365
transform -1 0 42784 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_4  _1028_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1029_
timestamp 1698431365
transform -1 0 42336 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  _1030_
timestamp 1698431365
transform 1 0 42112 0 1 23520
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1031_
timestamp 1698431365
transform 1 0 42448 0 -1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1032_
timestamp 1698431365
transform -1 0 46480 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1033_
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1034_
timestamp 1698431365
transform -1 0 52304 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1035_
timestamp 1698431365
transform 1 0 50848 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1036_
timestamp 1698431365
transform 1 0 44240 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1037_
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1038_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 50176 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1039_
timestamp 1698431365
transform -1 0 29232 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1040_
timestamp 1698431365
transform 1 0 47152 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1041_
timestamp 1698431365
transform 1 0 47600 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1042_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1043_
timestamp 1698431365
transform 1 0 45248 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1044_
timestamp 1698431365
transform -1 0 45248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1045_
timestamp 1698431365
transform 1 0 45472 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1046_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1047_
timestamp 1698431365
transform 1 0 31024 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1048_
timestamp 1698431365
transform 1 0 38528 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1049_
timestamp 1698431365
transform 1 0 25312 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1050_
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1051_
timestamp 1698431365
transform -1 0 26656 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1052_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 -1 20384
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1053_
timestamp 1698431365
transform 1 0 39536 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1054_
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1055_
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1056_
timestamp 1698431365
transform 1 0 38976 0 1 7840
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1057_
timestamp 1698431365
transform 1 0 45136 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1058_
timestamp 1698431365
transform -1 0 45696 0 1 3136
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1059_
timestamp 1698431365
transform 1 0 41104 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1060_
timestamp 1698431365
transform -1 0 45696 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1061_
timestamp 1698431365
transform -1 0 44240 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1062_
timestamp 1698431365
transform 1 0 39088 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1063_
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1064_
timestamp 1698431365
transform -1 0 41888 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1065_
timestamp 1698431365
transform 1 0 41776 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1066_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1067_
timestamp 1698431365
transform 1 0 41776 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1068_
timestamp 1698431365
transform -1 0 45920 0 -1 4704
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1069_
timestamp 1698431365
transform -1 0 39648 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1070_
timestamp 1698431365
transform 1 0 39648 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1071_
timestamp 1698431365
transform 1 0 42000 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1072_
timestamp 1698431365
transform -1 0 43120 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1073_
timestamp 1698431365
transform 1 0 38752 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1074_
timestamp 1698431365
transform -1 0 44464 0 1 4704
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1075_
timestamp 1698431365
transform -1 0 41776 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1076_
timestamp 1698431365
transform 1 0 37184 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1077_
timestamp 1698431365
transform -1 0 41888 0 1 6272
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1078_
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1079_
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1080_
timestamp 1698431365
transform 1 0 36960 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1081_
timestamp 1698431365
transform 1 0 37072 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1082_
timestamp 1698431365
transform -1 0 38752 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1083_
timestamp 1698431365
transform 1 0 36288 0 1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1084_
timestamp 1698431365
transform 1 0 36064 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1085_
timestamp 1698431365
transform -1 0 44912 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1086_
timestamp 1698431365
transform 1 0 47600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1087_
timestamp 1698431365
transform -1 0 4704 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1088_
timestamp 1698431365
transform -1 0 6272 0 -1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1089_
timestamp 1698431365
transform 1 0 49056 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1090_
timestamp 1698431365
transform 1 0 50400 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1091_
timestamp 1698431365
transform 1 0 8064 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1092_
timestamp 1698431365
transform 1 0 6160 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1093_
timestamp 1698431365
transform 1 0 50624 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1094_
timestamp 1698431365
transform -1 0 10416 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1095_
timestamp 1698431365
transform 1 0 50960 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1096_
timestamp 1698431365
transform -1 0 3696 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1097_
timestamp 1698431365
transform -1 0 6720 0 -1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1098_
timestamp 1698431365
transform 1 0 49952 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1099_
timestamp 1698431365
transform 1 0 50848 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1100_
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1101_
timestamp 1698431365
transform -1 0 58240 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1102_
timestamp 1698431365
transform -1 0 48944 0 1 4704
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1103_
timestamp 1698431365
transform -1 0 50176 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1104_
timestamp 1698431365
transform 1 0 45696 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1105_
timestamp 1698431365
transform 1 0 50400 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1106_
timestamp 1698431365
transform 1 0 50400 0 1 6272
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1107_
timestamp 1698431365
transform 1 0 51968 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1108_
timestamp 1698431365
transform -1 0 58352 0 1 4704
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1109_
timestamp 1698431365
transform 1 0 51184 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1110_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1111_
timestamp 1698431365
transform 1 0 52304 0 -1 9408
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1112_
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1113_
timestamp 1698431365
transform 1 0 56448 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1114_
timestamp 1698431365
transform -1 0 56224 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1115_
timestamp 1698431365
transform -1 0 58128 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1116_
timestamp 1698431365
transform 1 0 55104 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1117_
timestamp 1698431365
transform 1 0 53536 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1118_
timestamp 1698431365
transform 1 0 52976 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1119_
timestamp 1698431365
transform -1 0 58016 0 1 6272
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1120_
timestamp 1698431365
transform -1 0 58352 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1121_
timestamp 1698431365
transform -1 0 58128 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1122_
timestamp 1698431365
transform 1 0 56112 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1123_
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1124_
timestamp 1698431365
transform 1 0 54208 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1125_
timestamp 1698431365
transform -1 0 49840 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48832 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1127_
timestamp 1698431365
transform 1 0 47152 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1128_
timestamp 1698431365
transform -1 0 19824 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1129_
timestamp 1698431365
transform -1 0 10976 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1130_
timestamp 1698431365
transform -1 0 9968 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1131_
timestamp 1698431365
transform -1 0 10080 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1132_
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1133_
timestamp 1698431365
transform 1 0 10080 0 1 7840
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1134_
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1135_
timestamp 1698431365
transform -1 0 7616 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1136_
timestamp 1698431365
transform -1 0 4704 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1137_
timestamp 1698431365
transform -1 0 6608 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1138_
timestamp 1698431365
transform 1 0 5824 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1139_
timestamp 1698431365
transform 1 0 7616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1140_
timestamp 1698431365
transform 1 0 10304 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1141_
timestamp 1698431365
transform -1 0 14000 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1142_
timestamp 1698431365
transform 1 0 10080 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1143_
timestamp 1698431365
transform -1 0 14336 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1144_
timestamp 1698431365
transform 1 0 11760 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1145_
timestamp 1698431365
transform 1 0 12432 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1146_
timestamp 1698431365
transform -1 0 14336 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1147_
timestamp 1698431365
transform -1 0 8400 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1148_
timestamp 1698431365
transform -1 0 7616 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1149_
timestamp 1698431365
transform 1 0 2240 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1150_
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1151_
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1152_
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1153_
timestamp 1698431365
transform 1 0 5936 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1154_
timestamp 1698431365
transform -1 0 10080 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1155_
timestamp 1698431365
transform -1 0 12544 0 1 4704
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1156_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1157_
timestamp 1698431365
transform 1 0 3248 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1158_
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1159_
timestamp 1698431365
transform 1 0 4256 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1160_
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1161_
timestamp 1698431365
transform 1 0 3248 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1162_
timestamp 1698431365
transform 1 0 4592 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1163_
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1164_
timestamp 1698431365
transform -1 0 21168 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1165_
timestamp 1698431365
transform 1 0 21840 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1166_
timestamp 1698431365
transform -1 0 7056 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1167_
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1168_
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1169_
timestamp 1698431365
transform 1 0 7616 0 1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1170_
timestamp 1698431365
transform -1 0 9856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1171_
timestamp 1698431365
transform -1 0 9744 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1172_
timestamp 1698431365
transform -1 0 9072 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1173_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1174_
timestamp 1698431365
transform 1 0 22512 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1175_
timestamp 1698431365
transform -1 0 23744 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1176_
timestamp 1698431365
transform 1 0 22848 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1177_
timestamp 1698431365
transform 1 0 23184 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1178_
timestamp 1698431365
transform 1 0 21504 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1179_
timestamp 1698431365
transform 1 0 22064 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1180_
timestamp 1698431365
transform -1 0 26208 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1181_
timestamp 1698431365
transform 1 0 24304 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1182_
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1183_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1184_
timestamp 1698431365
transform -1 0 26880 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26208 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1186_
timestamp 1698431365
transform -1 0 25312 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1187_
timestamp 1698431365
transform -1 0 22736 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1188_
timestamp 1698431365
transform 1 0 22736 0 1 4704
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1189_
timestamp 1698431365
transform 1 0 14000 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1190_
timestamp 1698431365
transform 1 0 13552 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1191_
timestamp 1698431365
transform 1 0 14336 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1192_
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1193_
timestamp 1698431365
transform 1 0 14896 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1194_
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1195_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1196_
timestamp 1698431365
transform 1 0 13552 0 -1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1197_
timestamp 1698431365
transform 1 0 15344 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1198_
timestamp 1698431365
transform 1 0 12544 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1199_
timestamp 1698431365
transform -1 0 13664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1200_
timestamp 1698431365
transform 1 0 13104 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1201_
timestamp 1698431365
transform -1 0 10864 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1202_
timestamp 1698431365
transform 1 0 11760 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1203_
timestamp 1698431365
transform 1 0 6160 0 1 3136
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1204_
timestamp 1698431365
transform 1 0 7952 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1205_
timestamp 1698431365
transform -1 0 8848 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1206_
timestamp 1698431365
transform 1 0 7056 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1207_
timestamp 1698431365
transform -1 0 17024 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1208_
timestamp 1698431365
transform 1 0 23632 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1209_
timestamp 1698431365
transform -1 0 24752 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1210_
timestamp 1698431365
transform -1 0 19376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1211_
timestamp 1698431365
transform -1 0 5376 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1212_
timestamp 1698431365
transform -1 0 4256 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1213_
timestamp 1698431365
transform 1 0 4256 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1214_
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1215_
timestamp 1698431365
transform -1 0 22176 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1216_
timestamp 1698431365
transform 1 0 14000 0 -1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1217_
timestamp 1698431365
transform -1 0 19376 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1218_
timestamp 1698431365
transform 1 0 21504 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1219_
timestamp 1698431365
transform -1 0 19264 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1220_
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1221_
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1222_
timestamp 1698431365
transform 1 0 17808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1223_
timestamp 1698431365
transform -1 0 19600 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1224_
timestamp 1698431365
transform 1 0 18816 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1225_
timestamp 1698431365
transform -1 0 20272 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1226_
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1227_
timestamp 1698431365
transform -1 0 23296 0 -1 4704
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1228_
timestamp 1698431365
transform 1 0 20496 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1229_
timestamp 1698431365
transform 1 0 23296 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1230_
timestamp 1698431365
transform 1 0 26320 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1231_
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1232_
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1233_
timestamp 1698431365
transform -1 0 25984 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1234_
timestamp 1698431365
transform 1 0 26992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1235_
timestamp 1698431365
transform -1 0 27552 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1236_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1237_
timestamp 1698431365
transform 1 0 19936 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1238_
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1239_
timestamp 1698431365
transform 1 0 30464 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1240_
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1241_
timestamp 1698431365
transform -1 0 33152 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1242_
timestamp 1698431365
transform 1 0 31360 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1243_
timestamp 1698431365
transform 1 0 30352 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1244_
timestamp 1698431365
transform -1 0 28336 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1245_
timestamp 1698431365
transform -1 0 27664 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1246_
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1247_
timestamp 1698431365
transform -1 0 29904 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1248_
timestamp 1698431365
transform 1 0 29680 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1249_
timestamp 1698431365
transform -1 0 28672 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1250_
timestamp 1698431365
transform 1 0 30912 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1251_
timestamp 1698431365
transform 1 0 31584 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1252_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1253_
timestamp 1698431365
transform 1 0 34272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1254_
timestamp 1698431365
transform 1 0 33488 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1255_
timestamp 1698431365
transform 1 0 32368 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1256_
timestamp 1698431365
transform 1 0 31472 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1257_
timestamp 1698431365
transform 1 0 32592 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1258_
timestamp 1698431365
transform 1 0 33824 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1259_
timestamp 1698431365
transform 1 0 34720 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1260_
timestamp 1698431365
transform -1 0 31024 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1261_
timestamp 1698431365
transform 1 0 50960 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1262_
timestamp 1698431365
transform 1 0 49280 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1263_
timestamp 1698431365
transform 1 0 51296 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1264_
timestamp 1698431365
transform 1 0 52192 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1265_
timestamp 1698431365
transform 1 0 51856 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1266_
timestamp 1698431365
transform 1 0 53088 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1267_
timestamp 1698431365
transform 1 0 54320 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1268_
timestamp 1698431365
transform -1 0 56784 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1269_
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1270_
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1271_
timestamp 1698431365
transform 1 0 42672 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1272_
timestamp 1698431365
transform 1 0 44240 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1273_
timestamp 1698431365
transform 1 0 41888 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1274_
timestamp 1698431365
transform 1 0 47376 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1275_
timestamp 1698431365
transform 1 0 46480 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and4_4  _1276_
timestamp 1698431365
transform 1 0 49504 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1277_
timestamp 1698431365
transform 1 0 49056 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1278_
timestamp 1698431365
transform 1 0 42336 0 -1 23520
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1279_
timestamp 1698431365
transform -1 0 48272 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1280_
timestamp 1698431365
transform -1 0 50624 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1281_
timestamp 1698431365
transform -1 0 51296 0 1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1282_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1283_
timestamp 1698431365
transform -1 0 48384 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _1284_
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1285_
timestamp 1698431365
transform 1 0 43232 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1286_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42448 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1287_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 -1 18816
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1288_
timestamp 1698431365
transform 1 0 42000 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1289_
timestamp 1698431365
transform -1 0 43456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1290_
timestamp 1698431365
transform 1 0 42112 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1291_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42336 0 -1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1292_
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1293_
timestamp 1698431365
transform -1 0 52640 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1294_
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1295_
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1296_
timestamp 1698431365
transform -1 0 51968 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1297_
timestamp 1698431365
transform -1 0 48384 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1298_
timestamp 1698431365
transform 1 0 46144 0 1 17248
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1299_
timestamp 1698431365
transform 1 0 52640 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1300_
timestamp 1698431365
transform -1 0 48384 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1301_
timestamp 1698431365
transform 1 0 44912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1302_
timestamp 1698431365
transform -1 0 53088 0 -1 18816
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1303_
timestamp 1698431365
transform 1 0 48384 0 1 15680
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1304_
timestamp 1698431365
transform 1 0 51184 0 -1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1305_
timestamp 1698431365
transform 1 0 51968 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1306_
timestamp 1698431365
transform 1 0 53088 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1307_
timestamp 1698431365
transform 1 0 54432 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1308_
timestamp 1698431365
transform 1 0 54208 0 1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1309_
timestamp 1698431365
transform 1 0 51744 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1310_
timestamp 1698431365
transform 1 0 55440 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1311_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 54880 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1312_
timestamp 1698431365
transform 1 0 56560 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1313_
timestamp 1698431365
transform 1 0 56896 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1314_
timestamp 1698431365
transform -1 0 58352 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _1315_
timestamp 1698431365
transform 1 0 53312 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1316_
timestamp 1698431365
transform 1 0 53648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1317_
timestamp 1698431365
transform 1 0 53536 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1318_
timestamp 1698431365
transform 1 0 53536 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1319_
timestamp 1698431365
transform 1 0 53312 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1320_
timestamp 1698431365
transform 1 0 55440 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1321_
timestamp 1698431365
transform 1 0 50848 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1322_
timestamp 1698431365
transform 1 0 53088 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1323_
timestamp 1698431365
transform -1 0 53424 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1324_
timestamp 1698431365
transform -1 0 54208 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1325_
timestamp 1698431365
transform 1 0 54992 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1326_
timestamp 1698431365
transform 1 0 53312 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1327_
timestamp 1698431365
transform -1 0 56112 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1328_
timestamp 1698431365
transform 1 0 55328 0 1 15680
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1329_
timestamp 1698431365
transform -1 0 58352 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1330_
timestamp 1698431365
transform 1 0 54208 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1331_
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1332_
timestamp 1698431365
transform 1 0 54768 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1333_
timestamp 1698431365
transform -1 0 58352 0 1 14112
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1334_
timestamp 1698431365
transform 1 0 47712 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1335_
timestamp 1698431365
transform -1 0 49952 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1336_
timestamp 1698431365
transform -1 0 49392 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1337_
timestamp 1698431365
transform -1 0 49840 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1338_
timestamp 1698431365
transform 1 0 48944 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1339_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 53424 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1340_
timestamp 1698431365
transform -1 0 7616 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1341_
timestamp 1698431365
transform 1 0 55104 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1342_
timestamp 1698431365
transform -1 0 56000 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1343_
timestamp 1698431365
transform -1 0 55104 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1344_
timestamp 1698431365
transform 1 0 34832 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1345_
timestamp 1698431365
transform 1 0 34832 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1346_
timestamp 1698431365
transform -1 0 51856 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1347_
timestamp 1698431365
transform -1 0 58352 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1348_
timestamp 1698431365
transform 1 0 54768 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1349_
timestamp 1698431365
transform 1 0 57232 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1350_
timestamp 1698431365
transform -1 0 56896 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1351_
timestamp 1698431365
transform 1 0 33264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1352_
timestamp 1698431365
transform -1 0 51744 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1353_
timestamp 1698431365
transform -1 0 58352 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1354_
timestamp 1698431365
transform 1 0 56896 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1355_
timestamp 1698431365
transform -1 0 56224 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1356_
timestamp 1698431365
transform 1 0 35392 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1357_
timestamp 1698431365
transform 1 0 50848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1358_
timestamp 1698431365
transform 1 0 55440 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1359_
timestamp 1698431365
transform -1 0 57568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1360_
timestamp 1698431365
transform -1 0 53648 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1361_
timestamp 1698431365
transform -1 0 36064 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1362_
timestamp 1698431365
transform 1 0 34832 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1363_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 53760 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1364_
timestamp 1698431365
transform 1 0 57792 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1365_
timestamp 1698431365
transform -1 0 29680 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1366_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1367_
timestamp 1698431365
transform 1 0 28224 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1368_
timestamp 1698431365
transform -1 0 47040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1369_
timestamp 1698431365
transform -1 0 42784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1370_
timestamp 1698431365
transform 1 0 42224 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1371_
timestamp 1698431365
transform 1 0 44912 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1372_
timestamp 1698431365
transform 1 0 45584 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1373_
timestamp 1698431365
transform 1 0 45696 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1374_
timestamp 1698431365
transform 1 0 47264 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1375_
timestamp 1698431365
transform 1 0 41104 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1376_
timestamp 1698431365
transform 1 0 41104 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1377_
timestamp 1698431365
transform 1 0 43568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1378_
timestamp 1698431365
transform 1 0 45584 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1379_
timestamp 1698431365
transform 1 0 47376 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1380_
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1381_
timestamp 1698431365
transform 1 0 49056 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1382_
timestamp 1698431365
transform 1 0 27888 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1383_
timestamp 1698431365
transform 1 0 26992 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1384_
timestamp 1698431365
transform 1 0 43792 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1385_
timestamp 1698431365
transform 1 0 46144 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1386_
timestamp 1698431365
transform 1 0 46704 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1387_
timestamp 1698431365
transform 1 0 47488 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1388_
timestamp 1698431365
transform 1 0 46816 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1389_
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1390_
timestamp 1698431365
transform -1 0 49280 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1391_
timestamp 1698431365
transform -1 0 49728 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0693__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0694__I
timestamp 1698431365
transform 1 0 5712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0695__A2
timestamp 1698431365
transform 1 0 6160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0700__B2
timestamp 1698431365
transform -1 0 2352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A2
timestamp 1698431365
transform 1 0 4816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0703__A3
timestamp 1698431365
transform 1 0 13552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0712__I
timestamp 1698431365
transform -1 0 2016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0714__A2
timestamp 1698431365
transform 1 0 5824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0715__B
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0717__A1
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0720__A2
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0721__A2
timestamp 1698431365
transform 1 0 7168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0721__A3
timestamp 1698431365
transform 1 0 6720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0725__A2
timestamp 1698431365
transform -1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__A2
timestamp 1698431365
transform -1 0 3584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__A3
timestamp 1698431365
transform -1 0 4480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0731__A1
timestamp 1698431365
transform 1 0 8064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0731__A2
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0732__I0
timestamp 1698431365
transform 1 0 13664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0735__A2
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0736__A2
timestamp 1698431365
transform 1 0 11536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__A3
timestamp 1698431365
transform 1 0 3472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0745__A1
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0745__A2
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0746__A1
timestamp 1698431365
transform 1 0 19600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0746__A2
timestamp 1698431365
transform 1 0 17584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0757__A2
timestamp 1698431365
transform -1 0 5376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0759__A1
timestamp 1698431365
transform -1 0 10528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0759__A3
timestamp 1698431365
transform 1 0 10864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0764__A3
timestamp 1698431365
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A2
timestamp 1698431365
transform 1 0 11424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0767__A3
timestamp 1698431365
transform -1 0 6384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0771__A1
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0773__A2
timestamp 1698431365
transform 1 0 13552 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0773__A3
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__A1
timestamp 1698431365
transform 1 0 7392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__A2
timestamp 1698431365
transform 1 0 7840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__B
timestamp 1698431365
transform 1 0 9856 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A1
timestamp 1698431365
transform -1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__B
timestamp 1698431365
transform 1 0 10304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__A1
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__A2
timestamp 1698431365
transform -1 0 10864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__B
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0780__A1
timestamp 1698431365
transform -1 0 7168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0780__A2
timestamp 1698431365
transform -1 0 5936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0782__A1
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0782__A2
timestamp 1698431365
transform 1 0 9968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__A1
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__A2
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0784__A1
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0785__A1
timestamp 1698431365
transform -1 0 11312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0785__B
timestamp 1698431365
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__A2
timestamp 1698431365
transform 1 0 6048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0787__A1
timestamp 1698431365
transform -1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0787__A2
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0790__A2
timestamp 1698431365
transform 1 0 5824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0792__A1
timestamp 1698431365
transform 1 0 14112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0792__B
timestamp 1698431365
transform 1 0 14560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0795__A2
timestamp 1698431365
transform -1 0 11312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0796__I0
timestamp 1698431365
transform 1 0 15680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0797__A2
timestamp 1698431365
transform 1 0 23072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0801__A2
timestamp 1698431365
transform -1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0808__A1
timestamp 1698431365
transform -1 0 24192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0808__A2
timestamp 1698431365
transform 1 0 22064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__A1
timestamp 1698431365
transform 1 0 29568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__A2
timestamp 1698431365
transform 1 0 7168 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0817__A2
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__A1
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0822__I
timestamp 1698431365
transform 1 0 5264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A1
timestamp 1698431365
transform 1 0 15232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__B
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0831__I0
timestamp 1698431365
transform 1 0 18032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__A2
timestamp 1698431365
transform 1 0 10416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__A1
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__A2
timestamp 1698431365
transform -1 0 16464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__A1
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__A2
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__B
timestamp 1698431365
transform 1 0 11984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__I
timestamp 1698431365
transform 1 0 22512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__A1
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0853__B
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A3
timestamp 1698431365
transform -1 0 26096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A1
timestamp 1698431365
transform 1 0 34496 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__I
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__A1
timestamp 1698431365
transform 1 0 22960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__A1
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A1
timestamp 1698431365
transform 1 0 31024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__A1
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__B
timestamp 1698431365
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__A3
timestamp 1698431365
transform -1 0 26544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__A1
timestamp 1698431365
transform 1 0 27664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__B
timestamp 1698431365
transform 1 0 29344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A2
timestamp 1698431365
transform 1 0 31808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A1
timestamp 1698431365
transform 1 0 31024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A1
timestamp 1698431365
transform -1 0 25424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__S
timestamp 1698431365
transform 1 0 25424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0945__A1
timestamp 1698431365
transform 1 0 39312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0945__A2
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0946__A2
timestamp 1698431365
transform 1 0 39312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__A1
timestamp 1698431365
transform 1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__A1
timestamp 1698431365
transform 1 0 39760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0960__A2
timestamp 1698431365
transform 1 0 43456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__A1
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__A2
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A1
timestamp 1698431365
transform 1 0 26432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A2
timestamp 1698431365
transform 1 0 25872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__A3
timestamp 1698431365
transform -1 0 2352 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0970__A3
timestamp 1698431365
transform 1 0 7504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A2
timestamp 1698431365
transform 1 0 5712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A3
timestamp 1698431365
transform 1 0 5712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A1
timestamp 1698431365
transform 1 0 3136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__A1
timestamp 1698431365
transform 1 0 27328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__A2
timestamp 1698431365
transform -1 0 27104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__B
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__I
timestamp 1698431365
transform 1 0 46816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__A3
timestamp 1698431365
transform -1 0 47936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__A3
timestamp 1698431365
transform 1 0 5712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0978__A1
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A1
timestamp 1698431365
transform -1 0 27664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A2
timestamp 1698431365
transform -1 0 28112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__A1
timestamp 1698431365
transform 1 0 46256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__A2
timestamp 1698431365
transform -1 0 46032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__A1
timestamp 1698431365
transform 1 0 47488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__A2
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__B1
timestamp 1698431365
transform -1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__B2
timestamp 1698431365
transform 1 0 23744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0984__A3
timestamp 1698431365
transform 1 0 44352 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__A1
timestamp 1698431365
transform 1 0 18256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__A2
timestamp 1698431365
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A1
timestamp 1698431365
transform -1 0 25536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__B
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A2
timestamp 1698431365
transform 1 0 48048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A3
timestamp 1698431365
transform 1 0 47600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__A3
timestamp 1698431365
transform 1 0 30464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__S
timestamp 1698431365
transform 1 0 34720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0993__A2
timestamp 1698431365
transform 1 0 33600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0994__A1
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__A1
timestamp 1698431365
transform 1 0 35504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__A2
timestamp 1698431365
transform 1 0 35392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A2
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__A1
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__A2
timestamp 1698431365
transform 1 0 29232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__S
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A1
timestamp 1698431365
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A2
timestamp 1698431365
transform -1 0 41216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A3
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__A1
timestamp 1698431365
transform -1 0 43344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__A1
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A2
timestamp 1698431365
transform -1 0 45472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__A3
timestamp 1698431365
transform 1 0 51744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A1
timestamp 1698431365
transform 1 0 29456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A2
timestamp 1698431365
transform 1 0 26768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A1
timestamp 1698431365
transform 1 0 46928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A2
timestamp 1698431365
transform 1 0 46704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A1
timestamp 1698431365
transform -1 0 47600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1698431365
transform -1 0 25984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A2
timestamp 1698431365
transform 1 0 29232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__B1
timestamp 1698431365
transform 1 0 26208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__B2
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A2
timestamp 1698431365
transform -1 0 45248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A1
timestamp 1698431365
transform 1 0 44128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A1
timestamp 1698431365
transform -1 0 39088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A1
timestamp 1698431365
transform -1 0 39536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__B
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__B2
timestamp 1698431365
transform -1 0 41328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__B1
timestamp 1698431365
transform 1 0 36960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A2
timestamp 1698431365
transform 1 0 37632 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A2
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A1
timestamp 1698431365
transform 1 0 3920 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A2
timestamp 1698431365
transform 1 0 6272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__A2
timestamp 1698431365
transform 1 0 47376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A2
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A2
timestamp 1698431365
transform 1 0 6272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A2
timestamp 1698431365
transform 1 0 50400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A2
timestamp 1698431365
transform 1 0 6048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A2
timestamp 1698431365
transform -1 0 50400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__A2
timestamp 1698431365
transform -1 0 4592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__A2
timestamp 1698431365
transform -1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A2
timestamp 1698431365
transform 1 0 50064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A2
timestamp 1698431365
transform 1 0 51632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__B
timestamp 1698431365
transform 1 0 44912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A3
timestamp 1698431365
transform 1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__A2
timestamp 1698431365
transform -1 0 50400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A1
timestamp 1698431365
transform 1 0 52080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__A2
timestamp 1698431365
transform -1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__A1
timestamp 1698431365
transform 1 0 49952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform -1 0 47152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A2
timestamp 1698431365
transform 1 0 48832 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__B
timestamp 1698431365
transform 1 0 49056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__A1
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1698431365
transform 1 0 11200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1130__A2
timestamp 1698431365
transform 1 0 9968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__A1
timestamp 1698431365
transform -1 0 3696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__A2
timestamp 1698431365
transform -1 0 3248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__I0
timestamp 1698431365
transform -1 0 4144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A1
timestamp 1698431365
transform -1 0 6720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A1
timestamp 1698431365
transform 1 0 12544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__A1
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__A2
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__A1
timestamp 1698431365
transform 1 0 7504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A1
timestamp 1698431365
transform -1 0 3584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A2
timestamp 1698431365
transform -1 0 4032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__A1
timestamp 1698431365
transform 1 0 5600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A1
timestamp 1698431365
transform 1 0 5488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__A1
timestamp 1698431365
transform 1 0 3360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__A1
timestamp 1698431365
transform -1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A2
timestamp 1698431365
transform 1 0 21616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__A1
timestamp 1698431365
transform 1 0 6272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__A1
timestamp 1698431365
transform 1 0 20160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A1
timestamp 1698431365
transform 1 0 21616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1180__A2
timestamp 1698431365
transform 1 0 26880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1183__A1
timestamp 1698431365
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1183__A2
timestamp 1698431365
transform 1 0 26432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A2
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__B
timestamp 1698431365
transform 1 0 22512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__A1
timestamp 1698431365
transform 1 0 13776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__A2
timestamp 1698431365
transform 1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__A1
timestamp 1698431365
transform 1 0 14672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__B
timestamp 1698431365
transform 1 0 15568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__C
timestamp 1698431365
transform 1 0 14896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__A1
timestamp 1698431365
transform 1 0 7168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__A1
timestamp 1698431365
transform 1 0 7728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__A2
timestamp 1698431365
transform -1 0 4816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__B
timestamp 1698431365
transform 1 0 5040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__B2
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1215__A1
timestamp 1698431365
transform 1 0 22400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1235__A1
timestamp 1698431365
transform 1 0 27776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__C
timestamp 1698431365
transform 1 0 25312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1241__A1
timestamp 1698431365
transform 1 0 32256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1257__A1
timestamp 1698431365
transform 1 0 32368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A2
timestamp 1698431365
transform 1 0 31024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A1
timestamp 1698431365
transform 1 0 50736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A2
timestamp 1698431365
transform 1 0 49840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A3
timestamp 1698431365
transform 1 0 50288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A1
timestamp 1698431365
transform 1 0 50400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A2
timestamp 1698431365
transform 1 0 49504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__A2
timestamp 1698431365
transform 1 0 52976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__A2
timestamp 1698431365
transform 1 0 53424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__A2
timestamp 1698431365
transform 1 0 52864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__A1
timestamp 1698431365
transform 1 0 55888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__A2
timestamp 1698431365
transform 1 0 54768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__A2
timestamp 1698431365
transform 1 0 52080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__A1
timestamp 1698431365
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__B2
timestamp 1698431365
transform 1 0 45360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__I
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__A1
timestamp 1698431365
transform 1 0 42112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__A1
timestamp 1698431365
transform 1 0 49280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__B2
timestamp 1698431365
transform 1 0 48832 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__B
timestamp 1698431365
transform 1 0 47488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1304__A1
timestamp 1698431365
transform 1 0 50960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__A2
timestamp 1698431365
transform -1 0 53088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__A1
timestamp 1698431365
transform 1 0 51632 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__A2
timestamp 1698431365
transform 1 0 54768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__A1
timestamp 1698431365
transform 1 0 55216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__A1
timestamp 1698431365
transform 1 0 56672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1321__A1
timestamp 1698431365
transform 1 0 50624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1327__A1
timestamp 1698431365
transform -1 0 55328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1327__A2
timestamp 1698431365
transform 1 0 54544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__A1
timestamp 1698431365
transform 1 0 48048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A1
timestamp 1698431365
transform 1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A2
timestamp 1698431365
transform -1 0 48384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__B
timestamp 1698431365
transform 1 0 50064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__A2
timestamp 1698431365
transform 1 0 55888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__B
timestamp 1698431365
transform -1 0 54768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__A2
timestamp 1698431365
transform 1 0 53760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__B
timestamp 1698431365
transform 1 0 53984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__A2
timestamp 1698431365
transform 1 0 34608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__A1
timestamp 1698431365
transform 1 0 52528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__A2
timestamp 1698431365
transform 1 0 52080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A2
timestamp 1698431365
transform 1 0 54656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__B
timestamp 1698431365
transform 1 0 53536 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__B
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__A1
timestamp 1698431365
transform 1 0 50624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__A2
timestamp 1698431365
transform 1 0 51968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__B
timestamp 1698431365
transform 1 0 58128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__B
timestamp 1698431365
transform 1 0 54880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A1
timestamp 1698431365
transform 1 0 49952 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A2
timestamp 1698431365
transform -1 0 50624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__B
timestamp 1698431365
transform 1 0 55216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__A3
timestamp 1698431365
transform 1 0 52080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A1
timestamp 1698431365
transform 1 0 52976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__B1
timestamp 1698431365
transform 1 0 53984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__B2
timestamp 1698431365
transform 1 0 54432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1365__I
timestamp 1698431365
transform 1 0 29904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__B
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1369__A2
timestamp 1698431365
transform 1 0 41664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A1
timestamp 1698431365
transform -1 0 42672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1698431365
transform 1 0 40880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__A1
timestamp 1698431365
transform 1 0 50848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__A2
timestamp 1698431365
transform 1 0 50400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__B2
timestamp 1698431365
transform 1 0 51296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1382__A3
timestamp 1698431365
transform 1 0 28224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__A1
timestamp 1698431365
transform -1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__A2
timestamp 1698431365
transform -1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__B2
timestamp 1698431365
transform 1 0 48832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 4256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 4368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 6944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 8400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 1904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 1792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 4704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 7952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 7952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 6048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 30688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 52192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output27_I
timestamp 1698431365
transform 1 0 56560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_16 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_20
timestamp 1698431365
transform 1 0 3584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_24
timestamp 1698431365
transform 1 0 4032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_28
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_32
timestamp 1698431365
transform 1 0 4928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_40
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_42 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6048 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_50
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_54 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7392 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_62
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_66
timestamp 1698431365
transform 1 0 8736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_110 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_126
timestamp 1698431365
transform 1 0 15456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_134
timestamp 1698431365
transform 1 0 16352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_188
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_196
timestamp 1698431365
transform 1 0 23296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698431365
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_211
timestamp 1698431365
transform 1 0 24976 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_220
timestamp 1698431365
transform 1 0 25984 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698431365
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_284
timestamp 1698431365
transform 1 0 33152 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_300
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_304
timestamp 1698431365
transform 1 0 35392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_327
timestamp 1698431365
transform 1 0 37968 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_335
timestamp 1698431365
transform 1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_350
timestamp 1698431365
transform 1 0 40544 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_354
timestamp 1698431365
transform 1 0 40992 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_373
timestamp 1698431365
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_396
timestamp 1698431365
transform 1 0 45696 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_404
timestamp 1698431365
transform 1 0 46592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_436
timestamp 1698431365
transform 1 0 50176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_440
timestamp 1698431365
transform 1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_507
timestamp 1698431365
transform 1 0 58128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1698431365
transform 1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_12
timestamp 1698431365
transform 1 0 2688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_14
timestamp 1698431365
transform 1 0 2912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_17
timestamp 1698431365
transform 1 0 3248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_21
timestamp 1698431365
transform 1 0 3696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_25
timestamp 1698431365
transform 1 0 4144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_36
timestamp 1698431365
transform 1 0 5376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_40
timestamp 1698431365
transform 1 0 5824 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_49
timestamp 1698431365
transform 1 0 6832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_63
timestamp 1698431365
transform 1 0 8400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_67
timestamp 1698431365
transform 1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_78
timestamp 1698431365
transform 1 0 10080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_92
timestamp 1698431365
transform 1 0 11648 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_169
timestamp 1698431365
transform 1 0 20272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_222
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_237
timestamp 1698431365
transform 1 0 27888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_239
timestamp 1698431365
transform 1 0 28112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_248
timestamp 1698431365
transform 1 0 29120 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_256
timestamp 1698431365
transform 1 0 30016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_288
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_304
timestamp 1698431365
transform 1 0 35392 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_308
timestamp 1698431365
transform 1 0 35840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_325
timestamp 1698431365
transform 1 0 37744 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_329
timestamp 1698431365
transform 1 0 38192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_331
timestamp 1698431365
transform 1 0 38416 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_342
timestamp 1698431365
transform 1 0 39648 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_354
timestamp 1698431365
transform 1 0 40992 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_360
timestamp 1698431365
transform 1 0 41664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_398
timestamp 1698431365
transform 1 0 45920 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_406
timestamp 1698431365
transform 1 0 46816 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_410
timestamp 1698431365
transform 1 0 47264 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_450
timestamp 1698431365
transform 1 0 51744 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_496
timestamp 1698431365
transform 1 0 56896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_498
timestamp 1698431365
transform 1 0 57120 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_10
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_14
timestamp 1698431365
transform 1 0 2912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_55
timestamp 1698431365
transform 1 0 7504 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_116
timestamp 1698431365
transform 1 0 14336 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_124
timestamp 1698431365
transform 1 0 15232 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_140
timestamp 1698431365
transform 1 0 17024 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_162
timestamp 1698431365
transform 1 0 19488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_166
timestamp 1698431365
transform 1 0 19936 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_185
timestamp 1698431365
transform 1 0 22064 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_228
timestamp 1698431365
transform 1 0 26880 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_257
timestamp 1698431365
transform 1 0 30128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_271
timestamp 1698431365
transform 1 0 31696 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_287
timestamp 1698431365
transform 1 0 33488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_291
timestamp 1698431365
transform 1 0 33936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_293
timestamp 1698431365
transform 1 0 34160 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_310
timestamp 1698431365
transform 1 0 36064 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698431365
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_321
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_323
timestamp 1698431365
transform 1 0 37520 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_397
timestamp 1698431365
transform 1 0 45808 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_425
timestamp 1698431365
transform 1 0 48944 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_436
timestamp 1698431365
transform 1 0 50176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_440
timestamp 1698431365
transform 1 0 50624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_444
timestamp 1698431365
transform 1 0 51072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_448
timestamp 1698431365
transform 1 0 51520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1698431365
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698431365
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_473
timestamp 1698431365
transform 1 0 54320 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_6
timestamp 1698431365
transform 1 0 2016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_16
timestamp 1698431365
transform 1 0 3136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_20
timestamp 1698431365
transform 1 0 3584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_24
timestamp 1698431365
transform 1 0 4032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_28
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_31
timestamp 1698431365
transform 1 0 4816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_35
timestamp 1698431365
transform 1 0 5264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_39
timestamp 1698431365
transform 1 0 5712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_41
timestamp 1698431365
transform 1 0 5936 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_44
timestamp 1698431365
transform 1 0 6272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_48
timestamp 1698431365
transform 1 0 6720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_52
timestamp 1698431365
transform 1 0 7168 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_56
timestamp 1698431365
transform 1 0 7616 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_67
timestamp 1698431365
transform 1 0 8848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_76
timestamp 1698431365
transform 1 0 9856 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_85
timestamp 1698431365
transform 1 0 10864 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_117
timestamp 1698431365
transform 1 0 14448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_133
timestamp 1698431365
transform 1 0 16240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_163
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_171
timestamp 1698431365
transform 1 0 20496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_175
timestamp 1698431365
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_177
timestamp 1698431365
transform 1 0 21168 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_186
timestamp 1698431365
transform 1 0 22176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_190
timestamp 1698431365
transform 1 0 22624 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_216
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_224
timestamp 1698431365
transform 1 0 26432 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_234
timestamp 1698431365
transform 1 0 27552 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_238
timestamp 1698431365
transform 1 0 28000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_242
timestamp 1698431365
transform 1 0 28448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_244
timestamp 1698431365
transform 1 0 28672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_247
timestamp 1698431365
transform 1 0 29008 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_263
timestamp 1698431365
transform 1 0 30800 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_267
timestamp 1698431365
transform 1 0 31248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_269
timestamp 1698431365
transform 1 0 31472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_288
timestamp 1698431365
transform 1 0 33600 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_296
timestamp 1698431365
transform 1 0 34496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_298
timestamp 1698431365
transform 1 0 34720 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_307
timestamp 1698431365
transform 1 0 35728 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_315
timestamp 1698431365
transform 1 0 36624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_317
timestamp 1698431365
transform 1 0 36848 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_336
timestamp 1698431365
transform 1 0 38976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_340
timestamp 1698431365
transform 1 0 39424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_360
timestamp 1698431365
transform 1 0 41664 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_377
timestamp 1698431365
transform 1 0 43568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_393
timestamp 1698431365
transform 1 0 45360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_395
timestamp 1698431365
transform 1 0 45584 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_432
timestamp 1698431365
transform 1 0 49728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_447
timestamp 1698431365
transform 1 0 51408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_451
timestamp 1698431365
transform 1 0 51856 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_457
timestamp 1698431365
transform 1 0 52528 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_465
timestamp 1698431365
transform 1 0 53424 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_494
timestamp 1698431365
transform 1 0 56672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_24
timestamp 1698431365
transform 1 0 4032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_28
timestamp 1698431365
transform 1 0 4480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_32
timestamp 1698431365
transform 1 0 4928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_60
timestamp 1698431365
transform 1 0 8064 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_76
timestamp 1698431365
transform 1 0 9856 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_79
timestamp 1698431365
transform 1 0 10192 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_95
timestamp 1698431365
transform 1 0 11984 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_160
timestamp 1698431365
transform 1 0 19264 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_193
timestamp 1698431365
transform 1 0 22960 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_214
timestamp 1698431365
transform 1 0 25312 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_230
timestamp 1698431365
transform 1 0 27104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_232
timestamp 1698431365
transform 1 0 27328 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_263
timestamp 1698431365
transform 1 0 30800 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_271
timestamp 1698431365
transform 1 0 31696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_275
timestamp 1698431365
transform 1 0 32144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_284
timestamp 1698431365
transform 1 0 33152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_286
timestamp 1698431365
transform 1 0 33376 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_292
timestamp 1698431365
transform 1 0 34048 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_296
timestamp 1698431365
transform 1 0 34496 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_309
timestamp 1698431365
transform 1 0 35952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_313
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_362
timestamp 1698431365
transform 1 0 41888 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_378
timestamp 1698431365
transform 1 0 43680 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_433
timestamp 1698431365
transform 1 0 49840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_437
timestamp 1698431365
transform 1 0 50288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_462
timestamp 1698431365
transform 1 0 53088 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_470
timestamp 1698431365
transform 1 0 53984 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_506
timestamp 1698431365
transform 1 0 58016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_508
timestamp 1698431365
transform 1 0 58240 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_30
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_36
timestamp 1698431365
transform 1 0 5376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_53
timestamp 1698431365
transform 1 0 7280 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_57
timestamp 1698431365
transform 1 0 7728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_61
timestamp 1698431365
transform 1 0 8176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_65
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_77
timestamp 1698431365
transform 1 0 9968 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_90
timestamp 1698431365
transform 1 0 11424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_92
timestamp 1698431365
transform 1 0 11648 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_132
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_146
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_155
timestamp 1698431365
transform 1 0 18704 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_163
timestamp 1698431365
transform 1 0 19600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_165
timestamp 1698431365
transform 1 0 19824 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_178
timestamp 1698431365
transform 1 0 21280 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_194
timestamp 1698431365
transform 1 0 23072 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_202
timestamp 1698431365
transform 1 0 23968 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_222
timestamp 1698431365
transform 1 0 26208 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_230
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_248
timestamp 1698431365
transform 1 0 29120 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_252
timestamp 1698431365
transform 1 0 29568 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_265
timestamp 1698431365
transform 1 0 31024 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_273
timestamp 1698431365
transform 1 0 31920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_301
timestamp 1698431365
transform 1 0 35056 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_317
timestamp 1698431365
transform 1 0 36848 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_325
timestamp 1698431365
transform 1 0 37744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_329
timestamp 1698431365
transform 1 0 38192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_331
timestamp 1698431365
transform 1 0 38416 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_410
timestamp 1698431365
transform 1 0 47264 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_414
timestamp 1698431365
transform 1 0 47712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_426 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49056 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_27
timestamp 1698431365
transform 1 0 4368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_33
timestamp 1698431365
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_97
timestamp 1698431365
transform 1 0 12208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_116
timestamp 1698431365
transform 1 0 14336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_120
timestamp 1698431365
transform 1 0 14784 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_133
timestamp 1698431365
transform 1 0 16240 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_149
timestamp 1698431365
transform 1 0 18032 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_157
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_173
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_203
timestamp 1698431365
transform 1 0 24080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_222
timestamp 1698431365
transform 1 0 26208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_226
timestamp 1698431365
transform 1 0 26656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_293
timestamp 1698431365
transform 1 0 34160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_297
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_309
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_330
timestamp 1698431365
transform 1 0 38304 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_334
timestamp 1698431365
transform 1 0 38752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_408
timestamp 1698431365
transform 1 0 47040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_428
timestamp 1698431365
transform 1 0 49280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_450
timestamp 1698431365
transform 1 0 51744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_493
timestamp 1698431365
transform 1 0 56560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_507
timestamp 1698431365
transform 1 0 58128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_36
timestamp 1698431365
transform 1 0 5376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_38
timestamp 1698431365
transform 1 0 5600 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_41
timestamp 1698431365
transform 1 0 5936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_43
timestamp 1698431365
transform 1 0 6160 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_53
timestamp 1698431365
transform 1 0 7280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_57
timestamp 1698431365
transform 1 0 7728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_61
timestamp 1698431365
transform 1 0 8176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_63
timestamp 1698431365
transform 1 0 8400 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_86
timestamp 1698431365
transform 1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_90
timestamp 1698431365
transform 1 0 11424 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_106
timestamp 1698431365
transform 1 0 13216 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_109
timestamp 1698431365
transform 1 0 13552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_113
timestamp 1698431365
transform 1 0 14000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_115
timestamp 1698431365
transform 1 0 14224 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_125
timestamp 1698431365
transform 1 0 15344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_161
timestamp 1698431365
transform 1 0 19376 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_177
timestamp 1698431365
transform 1 0 21168 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_228
timestamp 1698431365
transform 1 0 26880 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_244
timestamp 1698431365
transform 1 0 28672 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_260
timestamp 1698431365
transform 1 0 30464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_264
timestamp 1698431365
transform 1 0 30912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_267
timestamp 1698431365
transform 1 0 31248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_275
timestamp 1698431365
transform 1 0 32144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_323
timestamp 1698431365
transform 1 0 37520 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_341
timestamp 1698431365
transform 1 0 39536 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698431365
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_365
timestamp 1698431365
transform 1 0 42224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_369
timestamp 1698431365
transform 1 0 42672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_403
timestamp 1698431365
transform 1 0 46480 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_409
timestamp 1698431365
transform 1 0 47152 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_428
timestamp 1698431365
transform 1 0 49280 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_436
timestamp 1698431365
transform 1 0 50176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_449
timestamp 1698431365
transform 1 0 51632 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_507
timestamp 1698431365
transform 1 0 58128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_16
timestamp 1698431365
transform 1 0 3136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_52
timestamp 1698431365
transform 1 0 7168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_63
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_65
timestamp 1698431365
transform 1 0 8624 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_75
timestamp 1698431365
transform 1 0 9744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_79
timestamp 1698431365
transform 1 0 10192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_83
timestamp 1698431365
transform 1 0 10640 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_89
timestamp 1698431365
transform 1 0 11312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_93
timestamp 1698431365
transform 1 0 11760 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_97
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_99
timestamp 1698431365
transform 1 0 12432 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_117
timestamp 1698431365
transform 1 0 14448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_134
timestamp 1698431365
transform 1 0 16352 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_142
timestamp 1698431365
transform 1 0 17248 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_146
timestamp 1698431365
transform 1 0 17696 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_149
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_169
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_226
timestamp 1698431365
transform 1 0 26656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_230
timestamp 1698431365
transform 1 0 27104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_232
timestamp 1698431365
transform 1 0 27328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_235
timestamp 1698431365
transform 1 0 27664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_239
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_255
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_283
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_285
timestamp 1698431365
transform 1 0 33264 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_374
timestamp 1698431365
transform 1 0 43232 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_378
timestamp 1698431365
transform 1 0 43680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_413
timestamp 1698431365
transform 1 0 47600 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_424
timestamp 1698431365
transform 1 0 48832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_432
timestamp 1698431365
transform 1 0 49728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_436
timestamp 1698431365
transform 1 0 50176 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_452
timestamp 1698431365
transform 1 0 51968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_465
timestamp 1698431365
transform 1 0 53424 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_469
timestamp 1698431365
transform 1 0 53872 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_471
timestamp 1698431365
transform 1 0 54096 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_6
timestamp 1698431365
transform 1 0 2016 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_122
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_156
timestamp 1698431365
transform 1 0 18816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_177
timestamp 1698431365
transform 1 0 21168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_179
timestamp 1698431365
transform 1 0 21392 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_200
timestamp 1698431365
transform 1 0 23744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_204
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_216
timestamp 1698431365
transform 1 0 25536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_230
timestamp 1698431365
transform 1 0 27104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_234
timestamp 1698431365
transform 1 0 27552 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_253
timestamp 1698431365
transform 1 0 29680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_257
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_259
timestamp 1698431365
transform 1 0 30352 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_262
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_266
timestamp 1698431365
transform 1 0 31136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_292
timestamp 1698431365
transform 1 0 34048 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_325
timestamp 1698431365
transform 1 0 37744 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_329
timestamp 1698431365
transform 1 0 38192 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_366
timestamp 1698431365
transform 1 0 42336 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_370
timestamp 1698431365
transform 1 0 42784 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_398
timestamp 1698431365
transform 1 0 45920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_400
timestamp 1698431365
transform 1 0 46144 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_407
timestamp 1698431365
transform 1 0 46928 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_426
timestamp 1698431365
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_436
timestamp 1698431365
transform 1 0 50176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_440
timestamp 1698431365
transform 1 0 50624 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_444
timestamp 1698431365
transform 1 0 51072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_474
timestamp 1698431365
transform 1 0 54432 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_478
timestamp 1698431365
transform 1 0 54880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_480
timestamp 1698431365
transform 1 0 55104 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_494
timestamp 1698431365
transform 1 0 56672 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_4
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_17
timestamp 1698431365
transform 1 0 3248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_21
timestamp 1698431365
transform 1 0 3696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_25
timestamp 1698431365
transform 1 0 4144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_29
timestamp 1698431365
transform 1 0 4592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_41
timestamp 1698431365
transform 1 0 5936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_80
timestamp 1698431365
transform 1 0 10304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_82
timestamp 1698431365
transform 1 0 10528 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_85
timestamp 1698431365
transform 1 0 10864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_95
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_113
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_116
timestamp 1698431365
transform 1 0 14336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_120
timestamp 1698431365
transform 1 0 14784 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_126
timestamp 1698431365
transform 1 0 15456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_130
timestamp 1698431365
transform 1 0 15904 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_146
timestamp 1698431365
transform 1 0 17696 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_154
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_156
timestamp 1698431365
transform 1 0 18816 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_165
timestamp 1698431365
transform 1 0 19824 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_191
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_197
timestamp 1698431365
transform 1 0 23408 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_220
timestamp 1698431365
transform 1 0 25984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_224
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_226
timestamp 1698431365
transform 1 0 26656 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1698431365
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_260
timestamp 1698431365
transform 1 0 30464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_262
timestamp 1698431365
transform 1 0 30688 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_286
timestamp 1698431365
transform 1 0 33376 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_302
timestamp 1698431365
transform 1 0 35168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_310
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_349
timestamp 1698431365
transform 1 0 40432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_353
timestamp 1698431365
transform 1 0 40880 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_374
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_399
timestamp 1698431365
transform 1 0 46032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_403
timestamp 1698431365
transform 1 0 46480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_410
timestamp 1698431365
transform 1 0 47264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_414
timestamp 1698431365
transform 1 0 47712 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_420
timestamp 1698431365
transform 1 0 48384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_424
timestamp 1698431365
transform 1 0 48832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_428
timestamp 1698431365
transform 1 0 49280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_432
timestamp 1698431365
transform 1 0 49728 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_438
timestamp 1698431365
transform 1 0 50400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_442
timestamp 1698431365
transform 1 0 50848 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_465
timestamp 1698431365
transform 1 0 53424 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_468
timestamp 1698431365
transform 1 0 53760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_472
timestamp 1698431365
transform 1 0 54208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_474
timestamp 1698431365
transform 1 0 54432 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_485
timestamp 1698431365
transform 1 0 55664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_507
timestamp 1698431365
transform 1 0 58128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_4
timestamp 1698431365
transform 1 0 1792 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_39
timestamp 1698431365
transform 1 0 5712 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_56
timestamp 1698431365
transform 1 0 7616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_62
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_76
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_92
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_107
timestamp 1698431365
transform 1 0 13328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_109
timestamp 1698431365
transform 1 0 13552 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_127
timestamp 1698431365
transform 1 0 15568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_131
timestamp 1698431365
transform 1 0 16016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_135
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_139
timestamp 1698431365
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_147
timestamp 1698431365
transform 1 0 17808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_161
timestamp 1698431365
transform 1 0 19376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_165
timestamp 1698431365
transform 1 0 19824 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_183
timestamp 1698431365
transform 1 0 21840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_187
timestamp 1698431365
transform 1 0 22288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_191
timestamp 1698431365
transform 1 0 22736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_205
timestamp 1698431365
transform 1 0 24304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_207
timestamp 1698431365
transform 1 0 24528 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_234
timestamp 1698431365
transform 1 0 27552 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_249
timestamp 1698431365
transform 1 0 29232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_253
timestamp 1698431365
transform 1 0 29680 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_261
timestamp 1698431365
transform 1 0 30576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_263
timestamp 1698431365
transform 1 0 30800 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_270
timestamp 1698431365
transform 1 0 31584 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_332
timestamp 1698431365
transform 1 0 38528 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_379
timestamp 1698431365
transform 1 0 43792 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_383
timestamp 1698431365
transform 1 0 44240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_396
timestamp 1698431365
transform 1 0 45696 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_404
timestamp 1698431365
transform 1 0 46592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_406
timestamp 1698431365
transform 1 0 46816 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_409
timestamp 1698431365
transform 1 0 47152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_433
timestamp 1698431365
transform 1 0 49840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_437
timestamp 1698431365
transform 1 0 50288 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_451
timestamp 1698431365
transform 1 0 51856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_455
timestamp 1698431365
transform 1 0 52304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_459
timestamp 1698431365
transform 1 0 52752 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_463
timestamp 1698431365
transform 1 0 53200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_467
timestamp 1698431365
transform 1 0 53648 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_470
timestamp 1698431365
transform 1 0 53984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_488
timestamp 1698431365
transform 1 0 56000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_16
timestamp 1698431365
transform 1 0 3136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_39
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_42
timestamp 1698431365
transform 1 0 6048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_46
timestamp 1698431365
transform 1 0 6496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_50
timestamp 1698431365
transform 1 0 6944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_54
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_74
timestamp 1698431365
transform 1 0 9632 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_78
timestamp 1698431365
transform 1 0 10080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_111
timestamp 1698431365
transform 1 0 13776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_117
timestamp 1698431365
transform 1 0 14448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_119
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_166
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_221
timestamp 1698431365
transform 1 0 26096 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_223
timestamp 1698431365
transform 1 0 26320 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_251
timestamp 1698431365
transform 1 0 29456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_259
timestamp 1698431365
transform 1 0 30352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_363
timestamp 1698431365
transform 1 0 42000 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_379
timestamp 1698431365
transform 1 0 43792 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_389
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_392
timestamp 1698431365
transform 1 0 45248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_401
timestamp 1698431365
transform 1 0 46256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_407
timestamp 1698431365
transform 1 0 46928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_415
timestamp 1698431365
transform 1 0 47824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_429
timestamp 1698431365
transform 1 0 49392 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_435
timestamp 1698431365
transform 1 0 50064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_439
timestamp 1698431365
transform 1 0 50512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_441
timestamp 1698431365
transform 1 0 50736 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_450
timestamp 1698431365
transform 1 0 51744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_454
timestamp 1698431365
transform 1 0 52192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_468
timestamp 1698431365
transform 1 0 53760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_472
timestamp 1698431365
transform 1 0 54208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_476
timestamp 1698431365
transform 1 0 54656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_51
timestamp 1698431365
transform 1 0 7056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_53
timestamp 1698431365
transform 1 0 7280 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_109
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_113
timestamp 1698431365
transform 1 0 14000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_115
timestamp 1698431365
transform 1 0 14224 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_148
timestamp 1698431365
transform 1 0 17920 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_152
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_191
timestamp 1698431365
transform 1 0 22736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_195
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_198
timestamp 1698431365
transform 1 0 23520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_202
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_218
timestamp 1698431365
transform 1 0 25760 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_231
timestamp 1698431365
transform 1 0 27216 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_233
timestamp 1698431365
transform 1 0 27440 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_247
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_251
timestamp 1698431365
transform 1 0 29456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_312
timestamp 1698431365
transform 1 0 36288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_373
timestamp 1698431365
transform 1 0 43120 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_381
timestamp 1698431365
transform 1 0 44016 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_398
timestamp 1698431365
transform 1 0 45920 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_414
timestamp 1698431365
transform 1 0 47712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_440
timestamp 1698431365
transform 1 0 50624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_442
timestamp 1698431365
transform 1 0 50848 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_469
timestamp 1698431365
transform 1 0 53872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_471
timestamp 1698431365
transform 1 0 54096 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_494
timestamp 1698431365
transform 1 0 56672 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_505
timestamp 1698431365
transform 1 0 57904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_15
timestamp 1698431365
transform 1 0 3024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_39
timestamp 1698431365
transform 1 0 5712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_42
timestamp 1698431365
transform 1 0 6048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_46
timestamp 1698431365
transform 1 0 6496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_48
timestamp 1698431365
transform 1 0 6720 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_75
timestamp 1698431365
transform 1 0 9744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_79
timestamp 1698431365
transform 1 0 10192 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_197
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_224
timestamp 1698431365
transform 1 0 26432 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_226
timestamp 1698431365
transform 1 0 26656 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_234
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_238
timestamp 1698431365
transform 1 0 28000 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_259
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_343
timestamp 1698431365
transform 1 0 39760 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_347
timestamp 1698431365
transform 1 0 40208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_368
timestamp 1698431365
transform 1 0 42560 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_429
timestamp 1698431365
transform 1 0 49392 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_433
timestamp 1698431365
transform 1 0 49840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_436
timestamp 1698431365
transform 1 0 50176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_440
timestamp 1698431365
transform 1 0 50624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_450
timestamp 1698431365
transform 1 0 51744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_452
timestamp 1698431365
transform 1 0 51968 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_467
timestamp 1698431365
transform 1 0 53648 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_471
timestamp 1698431365
transform 1 0 54096 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_45
timestamp 1698431365
transform 1 0 6384 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_51
timestamp 1698431365
transform 1 0 7056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_53
timestamp 1698431365
transform 1 0 7280 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_56
timestamp 1698431365
transform 1 0 7616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_144
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_199
timestamp 1698431365
transform 1 0 23632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_230
timestamp 1698431365
transform 1 0 27104 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_243
timestamp 1698431365
transform 1 0 28560 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_259
timestamp 1698431365
transform 1 0 30352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_261
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_286
timestamp 1698431365
transform 1 0 33376 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_309
timestamp 1698431365
transform 1 0 35952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_333
timestamp 1698431365
transform 1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_337
timestamp 1698431365
transform 1 0 39088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_341
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_370
timestamp 1698431365
transform 1 0 42784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_378
timestamp 1698431365
transform 1 0 43680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_382
timestamp 1698431365
transform 1 0 44128 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_390
timestamp 1698431365
transform 1 0 45024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_394
timestamp 1698431365
transform 1 0 45472 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_400
timestamp 1698431365
transform 1 0 46144 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_408
timestamp 1698431365
transform 1 0 47040 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_434
timestamp 1698431365
transform 1 0 49952 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_438
timestamp 1698431365
transform 1 0 50400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_454
timestamp 1698431365
transform 1 0 52192 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_462
timestamp 1698431365
transform 1 0 53088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_478
timestamp 1698431365
transform 1 0 54880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_482
timestamp 1698431365
transform 1 0 55328 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_488
timestamp 1698431365
transform 1 0 56000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_494
timestamp 1698431365
transform 1 0 56672 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_10
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_62
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_81
timestamp 1698431365
transform 1 0 10416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_189
timestamp 1698431365
transform 1 0 22512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_200
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_222
timestamp 1698431365
transform 1 0 26208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_260
timestamp 1698431365
transform 1 0 30464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_270
timestamp 1698431365
transform 1 0 31584 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_286
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_294
timestamp 1698431365
transform 1 0 34272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_303
timestamp 1698431365
transform 1 0 35280 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_358
timestamp 1698431365
transform 1 0 41440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_362
timestamp 1698431365
transform 1 0 41888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_370
timestamp 1698431365
transform 1 0 42784 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_374
timestamp 1698431365
transform 1 0 43232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_376
timestamp 1698431365
transform 1 0 43456 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_405
timestamp 1698431365
transform 1 0 46704 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_419
timestamp 1698431365
transform 1 0 48272 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_461
timestamp 1698431365
transform 1 0 52976 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_473
timestamp 1698431365
transform 1 0 54320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_4
timestamp 1698431365
transform 1 0 1792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_125
timestamp 1698431365
transform 1 0 15344 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_242
timestamp 1698431365
transform 1 0 28448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_246
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_304
timestamp 1698431365
transform 1 0 35392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_306
timestamp 1698431365
transform 1 0 35616 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_342
timestamp 1698431365
transform 1 0 39648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_344
timestamp 1698431365
transform 1 0 39872 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_362
timestamp 1698431365
transform 1 0 41888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_389
timestamp 1698431365
transform 1 0 44912 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_395
timestamp 1698431365
transform 1 0 45584 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_403
timestamp 1698431365
transform 1 0 46480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_426
timestamp 1698431365
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_430
timestamp 1698431365
transform 1 0 49504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_438
timestamp 1698431365
transform 1 0 50400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_442
timestamp 1698431365
transform 1 0 50848 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_489
timestamp 1698431365
transform 1 0 56112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_10
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_16
timestamp 1698431365
transform 1 0 3136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_23
timestamp 1698431365
transform 1 0 3920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_25
timestamp 1698431365
transform 1 0 4144 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_90
timestamp 1698431365
transform 1 0 11424 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_94
timestamp 1698431365
transform 1 0 11872 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_179
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_217
timestamp 1698431365
transform 1 0 25648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_263
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_291
timestamp 1698431365
transform 1 0 33936 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_321
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_340
timestamp 1698431365
transform 1 0 39424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_342
timestamp 1698431365
transform 1 0 39648 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_345
timestamp 1698431365
transform 1 0 39984 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_376
timestamp 1698431365
transform 1 0 43456 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_397
timestamp 1698431365
transform 1 0 45808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_399
timestamp 1698431365
transform 1 0 46032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_447
timestamp 1698431365
transform 1 0 51408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_4
timestamp 1698431365
transform 1 0 1792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_15
timestamp 1698431365
transform 1 0 3024 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_30
timestamp 1698431365
transform 1 0 4704 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_34
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_63
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_86
timestamp 1698431365
transform 1 0 10976 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_226
timestamp 1698431365
transform 1 0 26656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_250
timestamp 1698431365
transform 1 0 29344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_254
timestamp 1698431365
transform 1 0 29792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_271
timestamp 1698431365
transform 1 0 31696 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_293
timestamp 1698431365
transform 1 0 34160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_295
timestamp 1698431365
transform 1 0 34384 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_304
timestamp 1698431365
transform 1 0 35392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_341
timestamp 1698431365
transform 1 0 39536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_345
timestamp 1698431365
transform 1 0 39984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_347
timestamp 1698431365
transform 1 0 40208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_354
timestamp 1698431365
transform 1 0 40992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_462
timestamp 1698431365
transform 1 0 53088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_10
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_12
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_58
timestamp 1698431365
transform 1 0 7840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_170
timestamp 1698431365
transform 1 0 20384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698431365
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_454
timestamp 1698431365
transform 1 0 52192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_48
timestamp 1698431365
transform 1 0 6720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_263
timestamp 1698431365
transform 1 0 30800 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_333
timestamp 1698431365
transform 1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_337
timestamp 1698431365
transform 1 0 39088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_403
timestamp 1698431365
transform 1 0 46480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_432
timestamp 1698431365
transform 1 0 49728 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_476
timestamp 1698431365
transform 1 0 54656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_494
timestamp 1698431365
transform 1 0 56672 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_505
timestamp 1698431365
transform 1 0 57904 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_41
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_206
timestamp 1698431365
transform 1 0 24416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_226
timestamp 1698431365
transform 1 0 26656 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_256
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_263
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_267
timestamp 1698431365
transform 1 0 31248 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_271
timestamp 1698431365
transform 1 0 31696 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_304
timestamp 1698431365
transform 1 0 35392 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_475
timestamp 1698431365
transform 1 0 54544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_87
timestamp 1698431365
transform 1 0 11088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_89
timestamp 1698431365
transform 1 0 11312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_187
timestamp 1698431365
transform 1 0 22288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_263
timestamp 1698431365
transform 1 0 30800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_327
timestamp 1698431365
transform 1 0 37968 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_400
timestamp 1698431365
transform 1 0 46144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_402
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_479
timestamp 1698431365
transform 1 0 54992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_65
timestamp 1698431365
transform 1 0 8624 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_120
timestamp 1698431365
transform 1 0 14784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_162
timestamp 1698431365
transform 1 0 19488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_164
timestamp 1698431365
transform 1 0 19712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_211
timestamp 1698431365
transform 1 0 24976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_265
timestamp 1698431365
transform 1 0 31024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_267
timestamp 1698431365
transform 1 0 31248 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_292
timestamp 1698431365
transform 1 0 34048 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_308
timestamp 1698431365
transform 1 0 35840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_471
timestamp 1698431365
transform 1 0 54096 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_192
timestamp 1698431365
transform 1 0 22848 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_222
timestamp 1698431365
transform 1 0 26208 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_315
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_339
timestamp 1698431365
transform 1 0 39312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_341
timestamp 1698431365
transform 1 0 39536 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_388
timestamp 1698431365
transform 1 0 44800 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_392
timestamp 1698431365
transform 1 0 45248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_459
timestamp 1698431365
transform 1 0 52752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_463
timestamp 1698431365
transform 1 0 53200 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_472
timestamp 1698431365
transform 1 0 54208 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_485
timestamp 1698431365
transform 1 0 55664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_489
timestamp 1698431365
transform 1 0 56112 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_506
timestamp 1698431365
transform 1 0 58016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_6
timestamp 1698431365
transform 1 0 2016 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_111
timestamp 1698431365
transform 1 0 13776 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_227
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_229
timestamp 1698431365
transform 1 0 26992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_256
timestamp 1698431365
transform 1 0 30016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_286
timestamp 1698431365
transform 1 0 33376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_290
timestamp 1698431365
transform 1 0 33824 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_321
timestamp 1698431365
transform 1 0 37296 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_362
timestamp 1698431365
transform 1 0 41888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_395
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_399
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_440
timestamp 1698431365
transform 1 0 50624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_451
timestamp 1698431365
transform 1 0 51856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_475
timestamp 1698431365
transform 1 0 54544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_479
timestamp 1698431365
transform 1 0 54992 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_481
timestamp 1698431365
transform 1 0 55216 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_14
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_33
timestamp 1698431365
transform 1 0 5040 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_181
timestamp 1698431365
transform 1 0 21616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_183
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_224
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_293
timestamp 1698431365
transform 1 0 34160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_297
timestamp 1698431365
transform 1 0 34608 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_345
timestamp 1698431365
transform 1 0 39984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_380
timestamp 1698431365
transform 1 0 43904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_382
timestamp 1698431365
transform 1 0 44128 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_412
timestamp 1698431365
transform 1 0 47488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_424
timestamp 1698431365
transform 1 0 48832 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_463
timestamp 1698431365
transform 1 0 53200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_467
timestamp 1698431365
transform 1 0 53648 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_471
timestamp 1698431365
transform 1 0 54096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_473
timestamp 1698431365
transform 1 0 54320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_483
timestamp 1698431365
transform 1 0 55440 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_487
timestamp 1698431365
transform 1 0 55888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_489
timestamp 1698431365
transform 1 0 56112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_500
timestamp 1698431365
transform 1 0 57344 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698431365
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_39
timestamp 1698431365
transform 1 0 5712 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_42
timestamp 1698431365
transform 1 0 6048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_87
timestamp 1698431365
transform 1 0 11088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_131
timestamp 1698431365
transform 1 0 16016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_203
timestamp 1698431365
transform 1 0 24080 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_249
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_303
timestamp 1698431365
transform 1 0 35280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_352
timestamp 1698431365
transform 1 0 40768 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_356
timestamp 1698431365
transform 1 0 41216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_371
timestamp 1698431365
transform 1 0 42896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_375
timestamp 1698431365
transform 1 0 43344 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_419
timestamp 1698431365
transform 1 0 48272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_459
timestamp 1698431365
transform 1 0 52752 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_489
timestamp 1698431365
transform 1 0 56112 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_505
timestamp 1698431365
transform 1 0 57904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_28
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_104
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_125
timestamp 1698431365
transform 1 0 15344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_165
timestamp 1698431365
transform 1 0 19824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_169
timestamp 1698431365
transform 1 0 20272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_192
timestamp 1698431365
transform 1 0 22848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_210
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_214
timestamp 1698431365
transform 1 0 25312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_217
timestamp 1698431365
transform 1 0 25648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_221
timestamp 1698431365
transform 1 0 26096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_233
timestamp 1698431365
transform 1 0 27440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_237
timestamp 1698431365
transform 1 0 27888 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_248
timestamp 1698431365
transform 1 0 29120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_269
timestamp 1698431365
transform 1 0 31472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_271
timestamp 1698431365
transform 1 0 31696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_274
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_302
timestamp 1698431365
transform 1 0 35168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_334
timestamp 1698431365
transform 1 0 38752 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_338
timestamp 1698431365
transform 1 0 39200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_371
timestamp 1698431365
transform 1 0 42896 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_373
timestamp 1698431365
transform 1 0 43120 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_376
timestamp 1698431365
transform 1 0 43456 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_392
timestamp 1698431365
transform 1 0 45248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_400
timestamp 1698431365
transform 1 0 46144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_404
timestamp 1698431365
transform 1 0 46592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_410
timestamp 1698431365
transform 1 0 47264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_412
timestamp 1698431365
transform 1 0 47488 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_415
timestamp 1698431365
transform 1 0 47824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_448
timestamp 1698431365
transform 1 0 51520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_452
timestamp 1698431365
transform 1 0 51968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_456
timestamp 1698431365
transform 1 0 52416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_472
timestamp 1698431365
transform 1 0 54208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_478
timestamp 1698431365
transform 1 0 54880 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_490
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_505
timestamp 1698431365
transform 1 0 57904 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input4
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input5
timestamp 1698431365
transform -1 0 3136 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input6
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input7
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input8
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input11
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input12
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input13 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2688 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  input14
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  input15
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input16
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input17
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input18
timestamp 1698431365
transform 1 0 31248 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input19
timestamp 1698431365
transform 1 0 50176 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  load_slew28
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output20
timestamp 1698431365
transform 1 0 55328 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1698431365
transform 1 0 56784 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1698431365
transform 1 0 56784 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output23
timestamp 1698431365
transform -1 0 57904 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1698431365
transform 1 0 56784 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output25
timestamp 1698431365
transform 1 0 56784 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1698431365
transform -1 0 58352 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output27
timestamp 1698431365
transform 1 0 56784 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_30 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_31
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_32
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_33
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_34
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_35
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_36
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_37
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_38
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_39
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_40
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_41
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_42
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_43
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_44
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_45
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_46
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_47
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_48
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_49
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_50
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer1
timestamp 1698431365
transform 1 0 30352 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer2
timestamp 1698431365
transform 1 0 11312 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer3
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer4 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer5
timestamp 1698431365
transform -1 0 53536 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer6
timestamp 1698431365
transform -1 0 40544 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer7
timestamp 1698431365
transform 1 0 15456 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer8
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer9
timestamp 1698431365
transform -1 0 23296 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer10
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer11
timestamp 1698431365
transform -1 0 22512 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer12
timestamp 1698431365
transform -1 0 17920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer13
timestamp 1698431365
transform -1 0 16912 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer14
timestamp 1698431365
transform 1 0 23184 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer15
timestamp 1698431365
transform 1 0 39536 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  rebuffer16
timestamp 1698431365
transform 1 0 46144 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer17
timestamp 1698431365
transform -1 0 22288 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer18
timestamp 1698431365
transform 1 0 37856 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer19
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer20
timestamp 1698431365
transform 1 0 26544 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer21
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer22 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_60 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_61
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_62
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_63
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_64
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_65
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_66
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_67
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_68
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_69
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_70
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_71
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_72
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_73
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_74
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_75
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_76
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_77
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_78
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_79
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_80
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_81
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_82
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_83
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_84
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_85
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_86
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_87
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_88
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_89
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_90
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_91
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_92
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_93
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_94
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_95
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_96
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_97
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_98
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_99
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_100
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_101
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_102
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_103
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_104
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_105
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_106
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_107
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_108
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_109
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_110
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_111
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_112
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_113
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_114
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_115
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_116
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_117
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_118
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_119
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_120
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_121
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_122
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_123
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_124
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_125
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_126
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_127
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_128
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_129
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_130
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_131
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_132
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_133
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_134
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_135
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_137
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_138
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_139
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_144
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_149
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_150
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_154
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_155
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_156
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_157
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_158
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_159
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_160
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_161
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_162
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_163
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_164
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_165
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_166
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_167
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_168
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_169
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_170
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_171
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_172
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_173
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_174
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_175
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_176
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_177
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_178
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_179
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_180
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_181
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_182
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_183
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_184
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_185
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_186
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_187
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_188
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_189
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_190
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_193
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_194
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_195
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_198
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_199
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_200
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_206
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_209
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_210
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_211
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_212
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_213
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_214
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_215
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_216
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_217
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_218
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_219
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_220
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_221
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_222
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_223
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_224
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_225
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_226
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_227
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_228
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_229
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_230
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_231
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_232
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_233
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_234
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_235
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_236
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_237
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_238
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_239
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_240
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_241
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_242
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_243
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_244
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_245
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_246
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_247
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_248
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_249
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_250
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_251
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_252
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_253
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_254
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_255
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_256
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_257
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_258
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_259
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_260
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_261
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_262
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_263
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_264
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_265
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_266
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_267
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_268
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_269
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_270
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_271
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_272
timestamp 1698431365
transform 1 0 12768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_273
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_274
timestamp 1698431365
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_275
timestamp 1698431365
transform 1 0 24192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_276
timestamp 1698431365
transform 1 0 28000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_277
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_278
timestamp 1698431365
transform 1 0 35616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_279
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_280
timestamp 1698431365
transform 1 0 43232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_281
timestamp 1698431365
transform 1 0 47040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_282
timestamp 1698431365
transform 1 0 50848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_283
timestamp 1698431365
transform 1 0 54656 0 -1 26656
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 1344 800 1456 0 FreeSans 448 0 0 0 a[0]
port 0 nsew signal input
flabel metal3 s 0 3136 800 3248 0 FreeSans 448 0 0 0 a[1]
port 1 nsew signal input
flabel metal3 s 0 4928 800 5040 0 FreeSans 448 0 0 0 a[2]
port 2 nsew signal input
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 a[3]
port 3 nsew signal input
flabel metal3 s 0 8512 800 8624 0 FreeSans 448 0 0 0 a[4]
port 4 nsew signal input
flabel metal3 s 0 10304 800 10416 0 FreeSans 448 0 0 0 a[5]
port 5 nsew signal input
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 a[6]
port 6 nsew signal input
flabel metal3 s 0 13888 800 14000 0 FreeSans 448 0 0 0 a[7]
port 7 nsew signal input
flabel metal3 s 0 15680 800 15792 0 FreeSans 448 0 0 0 b[0]
port 8 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 b[1]
port 9 nsew signal input
flabel metal3 s 0 19264 800 19376 0 FreeSans 448 0 0 0 b[2]
port 10 nsew signal input
flabel metal3 s 0 21056 800 21168 0 FreeSans 448 0 0 0 b[3]
port 11 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 b[4]
port 12 nsew signal input
flabel metal3 s 0 24640 800 24752 0 FreeSans 448 0 0 0 b[5]
port 13 nsew signal input
flabel metal3 s 0 26432 800 26544 0 FreeSans 448 0 0 0 b[6]
port 14 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 b[7]
port 15 nsew signal input
flabel metal2 s 9856 29200 9968 30000 0 FreeSans 448 90 0 0 op[0]
port 16 nsew signal input
flabel metal2 s 29792 29200 29904 30000 0 FreeSans 448 90 0 0 op[1]
port 17 nsew signal input
flabel metal2 s 49728 29200 49840 30000 0 FreeSans 448 90 0 0 op[2]
port 18 nsew signal input
flabel metal3 s 59200 2240 60000 2352 0 FreeSans 448 0 0 0 out[0]
port 19 nsew signal tristate
flabel metal3 s 59200 5824 60000 5936 0 FreeSans 448 0 0 0 out[1]
port 20 nsew signal tristate
flabel metal3 s 59200 9408 60000 9520 0 FreeSans 448 0 0 0 out[2]
port 21 nsew signal tristate
flabel metal3 s 59200 12992 60000 13104 0 FreeSans 448 0 0 0 out[3]
port 22 nsew signal tristate
flabel metal3 s 59200 16576 60000 16688 0 FreeSans 448 0 0 0 out[4]
port 23 nsew signal tristate
flabel metal3 s 59200 20160 60000 20272 0 FreeSans 448 0 0 0 out[5]
port 24 nsew signal tristate
flabel metal3 s 59200 23744 60000 23856 0 FreeSans 448 0 0 0 out[6]
port 25 nsew signal tristate
flabel metal3 s 59200 27328 60000 27440 0 FreeSans 448 0 0 0 out[7]
port 26 nsew signal tristate
flabel metal4 s 8337 3076 8657 26716 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 22644 3076 22964 26716 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 36951 3076 37271 26716 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 51258 3076 51578 26716 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 15490 3076 15810 26716 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
flabel metal4 s 29797 3076 30117 26716 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
flabel metal4 s 44104 3076 44424 26716 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
flabel metal4 s 58411 3076 58731 26716 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 29960 25872 29960 25872 0 vdd
rlabel via1 30037 26656 30037 26656 0 vss
rlabel metal2 11032 20048 11032 20048 0 _0000_
rlabel metal2 13944 23072 13944 23072 0 _0001_
rlabel metal2 12040 22680 12040 22680 0 _0002_
rlabel metal2 12824 21280 12824 21280 0 _0003_
rlabel metal2 15624 19656 15624 19656 0 _0004_
rlabel metal2 25368 21448 25368 21448 0 _0005_
rlabel metal3 9912 19208 9912 19208 0 _0006_
rlabel metal2 12712 15624 12712 15624 0 _0007_
rlabel metal2 18088 15680 18088 15680 0 _0008_
rlabel metal2 15064 16352 15064 16352 0 _0009_
rlabel metal3 12040 15288 12040 15288 0 _0010_
rlabel metal2 14280 17192 14280 17192 0 _0011_
rlabel metal3 15680 19432 15680 19432 0 _0012_
rlabel metal3 13776 17080 13776 17080 0 _0013_
rlabel metal2 12712 17696 12712 17696 0 _0014_
rlabel metal3 13608 18536 13608 18536 0 _0015_
rlabel metal2 9128 18760 9128 18760 0 _0016_
rlabel metal2 14840 19320 14840 19320 0 _0017_
rlabel metal2 17528 12040 17528 12040 0 _0018_
rlabel metal2 10808 13440 10808 13440 0 _0019_
rlabel metal2 11144 14000 11144 14000 0 _0020_
rlabel metal3 11928 13048 11928 13048 0 _0021_
rlabel metal2 17080 12936 17080 12936 0 _0022_
rlabel metal2 12824 12992 12824 12992 0 _0023_
rlabel metal2 12488 13832 12488 13832 0 _0024_
rlabel metal2 15848 19992 15848 19992 0 _0025_
rlabel metal3 11704 21784 11704 21784 0 _0026_
rlabel metal2 20216 22904 20216 22904 0 _0027_
rlabel metal2 16576 19880 16576 19880 0 _0028_
rlabel metal2 20440 24528 20440 24528 0 _0029_
rlabel metal2 10808 9912 10808 9912 0 _0030_
rlabel metal2 13608 10920 13608 10920 0 _0031_
rlabel metal2 22680 23072 22680 23072 0 _0032_
rlabel metal3 21896 23352 21896 23352 0 _0033_
rlabel metal2 21672 24360 21672 24360 0 _0034_
rlabel metal2 26712 24192 26712 24192 0 _0035_
rlabel metal2 20888 23184 20888 23184 0 _0036_
rlabel metal2 26152 23576 26152 23576 0 _0037_
rlabel metal3 18592 26376 18592 26376 0 _0038_
rlabel metal2 26712 26432 26712 26432 0 _0039_
rlabel metal3 26488 22960 26488 22960 0 _0040_
rlabel metal2 26824 22848 26824 22848 0 _0041_
rlabel metal2 31416 22344 31416 22344 0 _0042_
rlabel metal2 35168 22568 35168 22568 0 _0043_
rlabel metal2 26376 19544 26376 19544 0 _0044_
rlabel metal2 24584 21448 24584 21448 0 _0045_
rlabel metal2 37576 17192 37576 17192 0 _0046_
rlabel metal2 21840 17528 21840 17528 0 _0047_
rlabel metal2 16632 20552 16632 20552 0 _0048_
rlabel metal2 16072 20720 16072 20720 0 _0049_
rlabel metal2 19320 18088 19320 18088 0 _0050_
rlabel metal3 9464 14728 9464 14728 0 _0051_
rlabel metal3 15372 16968 15372 16968 0 _0052_
rlabel metal3 16968 15176 16968 15176 0 _0053_
rlabel metal2 21112 13664 21112 13664 0 _0054_
rlabel metal2 18760 12936 18760 12936 0 _0055_
rlabel metal2 25256 15204 25256 15204 0 _0056_
rlabel metal2 18760 15400 18760 15400 0 _0057_
rlabel metal2 9576 17640 9576 17640 0 _0058_
rlabel metal2 17528 17696 17528 17696 0 _0059_
rlabel metal2 14616 22624 14616 22624 0 _0060_
rlabel metal2 17416 17304 17416 17304 0 _0061_
rlabel metal3 19992 16856 19992 16856 0 _0062_
rlabel metal2 23800 19488 23800 19488 0 _0063_
rlabel metal3 19376 13496 19376 13496 0 _0064_
rlabel metal2 22680 16072 22680 16072 0 _0065_
rlabel metal3 19040 16856 19040 16856 0 _0066_
rlabel metal2 23464 15204 23464 15204 0 _0067_
rlabel metal2 23128 16072 23128 16072 0 _0068_
rlabel metal3 22904 16968 22904 16968 0 _0069_
rlabel metal2 19432 19600 19432 19600 0 _0070_
rlabel metal2 17696 10584 17696 10584 0 _0071_
rlabel metal2 18648 16072 18648 16072 0 _0072_
rlabel metal2 17752 16968 17752 16968 0 _0073_
rlabel metal3 21056 18424 21056 18424 0 _0074_
rlabel metal2 21672 19768 21672 19768 0 _0075_
rlabel metal2 18200 20608 18200 20608 0 _0076_
rlabel metal2 22232 18592 22232 18592 0 _0077_
rlabel metal2 25592 17752 25592 17752 0 _0078_
rlabel metal2 19768 17640 19768 17640 0 _0079_
rlabel metal2 22792 14504 22792 14504 0 _0080_
rlabel metal3 23296 15176 23296 15176 0 _0081_
rlabel metal2 26152 16240 26152 16240 0 _0082_
rlabel metal2 33936 18424 33936 18424 0 _0083_
rlabel metal2 23464 16240 23464 16240 0 _0084_
rlabel metal2 35896 18704 35896 18704 0 _0085_
rlabel metal2 23408 13944 23408 13944 0 _0086_
rlabel metal2 23576 17024 23576 17024 0 _0087_
rlabel metal2 21560 17976 21560 17976 0 _0088_
rlabel metal2 37800 16408 37800 16408 0 _0089_
rlabel metal2 40152 13664 40152 13664 0 _0090_
rlabel metal2 23464 25480 23464 25480 0 _0091_
rlabel metal2 30184 23520 30184 23520 0 _0092_
rlabel metal2 26040 25984 26040 25984 0 _0093_
rlabel metal2 27832 24248 27832 24248 0 _0094_
rlabel metal2 36344 20160 36344 20160 0 _0095_
rlabel metal2 35112 19040 35112 19040 0 _0096_
rlabel metal3 26040 13720 26040 13720 0 _0097_
rlabel metal2 27664 12040 27664 12040 0 _0098_
rlabel metal2 26544 18536 26544 18536 0 _0099_
rlabel metal2 36232 19712 36232 19712 0 _0100_
rlabel metal2 39144 10864 39144 10864 0 _0101_
rlabel metal3 39088 12936 39088 12936 0 _0102_
rlabel metal2 26600 22064 26600 22064 0 _0103_
rlabel metal2 37016 21952 37016 21952 0 _0104_
rlabel metal2 24584 19544 24584 19544 0 _0105_
rlabel metal2 37576 20440 37576 20440 0 _0106_
rlabel metal2 37016 16184 37016 16184 0 _0107_
rlabel metal2 33768 24976 33768 24976 0 _0108_
rlabel metal2 25704 24024 25704 24024 0 _0109_
rlabel metal2 34832 15512 34832 15512 0 _0110_
rlabel metal2 34440 16184 34440 16184 0 _0111_
rlabel metal2 35784 13608 35784 13608 0 _0112_
rlabel metal2 35784 18480 35784 18480 0 _0113_
rlabel metal2 35224 15736 35224 15736 0 _0114_
rlabel metal2 35000 15568 35000 15568 0 _0115_
rlabel metal3 36960 13608 36960 13608 0 _0116_
rlabel metal2 35896 14728 35896 14728 0 _0117_
rlabel metal2 30856 21280 30856 21280 0 _0118_
rlabel metal2 32088 23800 32088 23800 0 _0119_
rlabel metal2 31416 17808 31416 17808 0 _0120_
rlabel metal2 30744 16856 30744 16856 0 _0121_
rlabel metal2 26488 17024 26488 17024 0 _0122_
rlabel metal2 30408 16240 30408 16240 0 _0123_
rlabel metal2 31192 16464 31192 16464 0 _0124_
rlabel metal2 31080 15568 31080 15568 0 _0125_
rlabel metal2 27384 23968 27384 23968 0 _0126_
rlabel metal3 27272 16072 27272 16072 0 _0127_
rlabel metal2 24808 19824 24808 19824 0 _0128_
rlabel metal2 27776 17080 27776 17080 0 _0129_
rlabel metal2 26264 17528 26264 17528 0 _0130_
rlabel metal3 25648 15848 25648 15848 0 _0131_
rlabel metal3 27048 16856 27048 16856 0 _0132_
rlabel metal2 27384 16016 27384 16016 0 _0133_
rlabel metal2 27720 15568 27720 15568 0 _0134_
rlabel metal2 28280 15232 28280 15232 0 _0135_
rlabel metal3 34664 14952 34664 14952 0 _0136_
rlabel metal2 32088 15568 32088 15568 0 _0137_
rlabel metal2 37016 15232 37016 15232 0 _0138_
rlabel metal3 39592 14392 39592 14392 0 _0139_
rlabel metal2 38248 15232 38248 15232 0 _0140_
rlabel metal2 38024 14336 38024 14336 0 _0141_
rlabel metal2 35112 12544 35112 12544 0 _0142_
rlabel metal2 32872 25424 32872 25424 0 _0143_
rlabel metal2 32760 25424 32760 25424 0 _0144_
rlabel metal2 31752 16520 31752 16520 0 _0145_
rlabel metal2 32872 17836 32872 17836 0 _0146_
rlabel metal3 29848 19208 29848 19208 0 _0147_
rlabel metal2 32704 19208 32704 19208 0 _0148_
rlabel metal3 31808 14504 31808 14504 0 _0149_
rlabel metal2 30744 14224 30744 14224 0 _0150_
rlabel metal3 33880 12152 33880 12152 0 _0151_
rlabel metal2 35896 12824 35896 12824 0 _0152_
rlabel metal2 36792 13048 36792 13048 0 _0153_
rlabel metal2 38696 14448 38696 14448 0 _0154_
rlabel metal2 41272 9016 41272 9016 0 _0155_
rlabel metal2 39144 11368 39144 11368 0 _0156_
rlabel metal2 39368 8456 39368 8456 0 _0157_
rlabel metal2 39144 6776 39144 6776 0 _0158_
rlabel metal2 30744 20272 30744 20272 0 _0159_
rlabel metal2 42392 19880 42392 19880 0 _0160_
rlabel metal3 33880 20664 33880 20664 0 _0161_
rlabel metal2 30520 19096 30520 19096 0 _0162_
rlabel metal2 39592 18928 39592 18928 0 _0163_
rlabel metal2 47992 19600 47992 19600 0 _0164_
rlabel metal3 24752 18424 24752 18424 0 _0165_
rlabel metal2 25928 18480 25928 18480 0 _0166_
rlabel metal2 25592 19264 25592 19264 0 _0167_
rlabel metal2 25144 20048 25144 20048 0 _0168_
rlabel metal2 22120 25032 22120 25032 0 _0169_
rlabel metal2 25256 25872 25256 25872 0 _0170_
rlabel metal3 25088 26152 25088 26152 0 _0171_
rlabel metal2 25032 22008 25032 22008 0 _0172_
rlabel metal2 26600 20384 26600 20384 0 _0173_
rlabel metal2 21560 21560 21560 21560 0 _0174_
rlabel metal2 22568 20720 22568 20720 0 _0175_
rlabel metal2 25368 19264 25368 19264 0 _0176_
rlabel metal2 22848 21560 22848 21560 0 _0177_
rlabel metal2 39032 15792 39032 15792 0 _0178_
rlabel metal2 23688 18312 23688 18312 0 _0179_
rlabel metal2 39256 16352 39256 16352 0 _0180_
rlabel metal2 40264 15680 40264 15680 0 _0181_
rlabel metal2 43288 24136 43288 24136 0 _0182_
rlabel metal2 35000 11256 35000 11256 0 _0183_
rlabel metal2 34888 11480 34888 11480 0 _0184_
rlabel metal2 31080 11256 31080 11256 0 _0185_
rlabel metal2 31192 11760 31192 11760 0 _0186_
rlabel metal2 39928 11144 39928 11144 0 _0187_
rlabel metal2 39760 11480 39760 11480 0 _0188_
rlabel metal2 36344 10920 36344 10920 0 _0189_
rlabel metal2 8904 16072 8904 16072 0 _0190_
rlabel metal2 40488 9856 40488 9856 0 _0191_
rlabel metal2 44072 21504 44072 21504 0 _0192_
rlabel metal2 41272 17136 41272 17136 0 _0193_
rlabel metal2 41048 17304 41048 17304 0 _0194_
rlabel metal2 42000 12040 42000 12040 0 _0195_
rlabel metal2 42952 10640 42952 10640 0 _0196_
rlabel metal2 46760 9464 46760 9464 0 _0197_
rlabel metal3 43512 9688 43512 9688 0 _0198_
rlabel metal2 43064 11312 43064 11312 0 _0199_
rlabel metal3 45920 9688 45920 9688 0 _0200_
rlabel metal2 12432 26264 12432 26264 0 _0201_
rlabel metal2 45192 10584 45192 10584 0 _0202_
rlabel metal3 41664 13496 41664 13496 0 _0203_
rlabel metal2 28392 14448 28392 14448 0 _0204_
rlabel metal3 34944 13720 34944 13720 0 _0205_
rlabel metal2 44744 11592 44744 11592 0 _0206_
rlabel metal2 7000 12768 7000 12768 0 _0207_
rlabel metal2 9128 10640 9128 10640 0 _0208_
rlabel metal2 2856 11088 2856 11088 0 _0209_
rlabel metal2 26488 13552 26488 13552 0 _0210_
rlabel metal3 26040 10584 26040 10584 0 _0211_
rlabel metal2 7784 24696 7784 24696 0 _0212_
rlabel metal2 44912 11480 44912 11480 0 _0213_
rlabel metal2 48776 26656 48776 26656 0 _0214_
rlabel metal2 49224 24752 49224 24752 0 _0215_
rlabel metal2 6664 10304 6664 10304 0 _0216_
rlabel metal2 4648 10304 4648 10304 0 _0217_
rlabel metal3 24696 10640 24696 10640 0 _0218_
rlabel metal2 47880 10640 47880 10640 0 _0219_
rlabel metal2 46760 10864 46760 10864 0 _0220_
rlabel metal2 47208 11200 47208 11200 0 _0221_
rlabel metal2 26768 13944 26768 13944 0 _0222_
rlabel metal2 9128 24584 9128 24584 0 _0223_
rlabel metal2 45640 12432 45640 12432 0 _0224_
rlabel metal2 26376 10136 26376 10136 0 _0225_
rlabel metal2 26600 10976 26600 10976 0 _0226_
rlabel metal2 50456 25816 50456 25816 0 _0227_
rlabel metal2 50232 22568 50232 22568 0 _0228_
rlabel metal3 41944 12656 41944 12656 0 _0229_
rlabel metal3 37016 23016 37016 23016 0 _0230_
rlabel metal2 39032 22624 39032 22624 0 _0231_
rlabel metal2 34104 25144 34104 25144 0 _0232_
rlabel metal2 33096 25424 33096 25424 0 _0233_
rlabel metal2 8904 24080 8904 24080 0 _0234_
rlabel metal2 41720 24360 41720 24360 0 _0235_
rlabel metal3 36624 18424 36624 18424 0 _0236_
rlabel metal3 38724 18424 38724 18424 0 _0237_
rlabel metal2 39368 23856 39368 23856 0 _0238_
rlabel metal2 39704 23688 39704 23688 0 _0239_
rlabel metal2 35784 24528 35784 24528 0 _0240_
rlabel metal2 38696 25200 38696 25200 0 _0241_
rlabel metal3 34384 23688 34384 23688 0 _0242_
rlabel metal2 35168 23800 35168 23800 0 _0243_
rlabel metal2 37576 24752 37576 24752 0 _0244_
rlabel metal2 2744 22624 2744 22624 0 _0245_
rlabel metal2 39144 20664 39144 20664 0 _0246_
rlabel metal2 35896 25144 35896 25144 0 _0247_
rlabel metal2 41048 22568 41048 22568 0 _0248_
rlabel metal2 40376 22792 40376 22792 0 _0249_
rlabel metal2 34552 20832 34552 20832 0 _0250_
rlabel metal2 44072 22176 44072 22176 0 _0251_
rlabel metal2 45976 22008 45976 22008 0 _0252_
rlabel metal2 28504 14168 28504 14168 0 _0253_
rlabel metal3 44576 14504 44576 14504 0 _0254_
rlabel metal2 37240 23128 37240 23128 0 _0255_
rlabel metal2 3752 23912 3752 23912 0 _0256_
rlabel metal2 46088 21504 46088 21504 0 _0257_
rlabel metal3 45360 19432 45360 19432 0 _0258_
rlabel metal2 46984 19936 46984 19936 0 _0259_
rlabel metal2 22792 21840 22792 21840 0 _0260_
rlabel metal2 23408 20104 23408 20104 0 _0261_
rlabel metal2 48776 18424 48776 18424 0 _0262_
rlabel metal2 43736 21224 43736 21224 0 _0263_
rlabel metal2 44744 25032 44744 25032 0 _0264_
rlabel metal2 44520 24976 44520 24976 0 _0265_
rlabel metal2 36008 25088 36008 25088 0 _0266_
rlabel metal2 4424 20496 4424 20496 0 _0267_
rlabel metal2 41384 25816 41384 25816 0 _0268_
rlabel metal2 43064 25368 43064 25368 0 _0269_
rlabel metal3 42616 24584 42616 24584 0 _0270_
rlabel metal3 44352 24696 44352 24696 0 _0271_
rlabel metal3 49672 23240 49672 23240 0 _0272_
rlabel metal3 42616 23128 42616 23128 0 _0273_
rlabel metal2 44744 21896 44744 21896 0 _0274_
rlabel metal2 45080 20720 45080 20720 0 _0275_
rlabel metal2 45080 18424 45080 18424 0 _0276_
rlabel metal3 52864 23240 52864 23240 0 _0277_
rlabel metal2 3192 24024 3192 24024 0 _0278_
rlabel metal2 51520 22568 51520 22568 0 _0279_
rlabel metal3 45024 15512 45024 15512 0 _0280_
rlabel metal2 44520 14728 44520 14728 0 _0281_
rlabel metal2 45024 13944 45024 13944 0 _0282_
rlabel metal2 50288 26040 50288 26040 0 _0283_
rlabel metal2 46760 13104 46760 13104 0 _0284_
rlabel metal2 47768 12656 47768 12656 0 _0285_
rlabel metal2 48048 12376 48048 12376 0 _0286_
rlabel metal2 45416 13384 45416 13384 0 _0287_
rlabel metal3 45080 13832 45080 13832 0 _0288_
rlabel metal2 16296 21840 16296 21840 0 _0289_
rlabel metal3 45248 12936 45248 12936 0 _0290_
rlabel metal2 40880 9240 40880 9240 0 _0291_
rlabel metal2 41944 4312 41944 4312 0 _0292_
rlabel metal2 39592 8624 39592 8624 0 _0293_
rlabel metal2 25592 22456 25592 22456 0 _0294_
rlabel metal2 24696 20664 24696 20664 0 _0295_
rlabel metal2 26152 18872 26152 18872 0 _0296_
rlabel metal2 40152 10696 40152 10696 0 _0297_
rlabel metal2 39816 10192 39816 10192 0 _0298_
rlabel metal2 16072 21952 16072 21952 0 _0299_
rlabel metal3 38864 9688 38864 9688 0 _0300_
rlabel metal2 41832 9072 41832 9072 0 _0301_
rlabel metal2 41216 4312 41216 4312 0 _0302_
rlabel metal2 46872 5488 46872 5488 0 _0303_
rlabel metal2 43624 5040 43624 5040 0 _0304_
rlabel metal3 42896 4312 42896 4312 0 _0305_
rlabel metal2 44744 7840 44744 7840 0 _0306_
rlabel metal2 43400 6664 43400 6664 0 _0307_
rlabel metal2 40600 14560 40600 14560 0 _0308_
rlabel metal2 41216 10696 41216 10696 0 _0309_
rlabel metal2 13608 26376 13608 26376 0 _0310_
rlabel metal2 41608 15232 41608 15232 0 _0311_
rlabel metal2 42280 9968 42280 9968 0 _0312_
rlabel metal2 43176 8512 43176 8512 0 _0313_
rlabel metal2 42672 4312 42672 4312 0 _0314_
rlabel metal3 45192 6664 45192 6664 0 _0315_
rlabel metal2 39480 5488 39480 5488 0 _0316_
rlabel metal2 40152 6384 40152 6384 0 _0317_
rlabel metal3 43568 6888 43568 6888 0 _0318_
rlabel metal2 42056 4368 42056 4368 0 _0319_
rlabel metal2 40040 4984 40040 4984 0 _0320_
rlabel metal2 5992 22680 5992 22680 0 _0321_
rlabel metal2 45864 6384 45864 6384 0 _0322_
rlabel metal2 40880 6664 40880 6664 0 _0323_
rlabel metal2 38248 6384 38248 6384 0 _0324_
rlabel metal2 45752 7000 45752 7000 0 _0325_
rlabel metal2 46984 7224 46984 7224 0 _0326_
rlabel metal3 41720 7560 41720 7560 0 _0327_
rlabel metal2 37296 8456 37296 8456 0 _0328_
rlabel metal2 37352 6384 37352 6384 0 _0329_
rlabel metal2 37856 3416 37856 3416 0 _0330_
rlabel metal2 36568 3920 36568 3920 0 _0331_
rlabel metal2 7672 25760 7672 25760 0 _0332_
rlabel metal3 39928 6720 39928 6720 0 _0333_
rlabel metal2 48776 6496 48776 6496 0 _0334_
rlabel metal2 49560 4256 49560 4256 0 _0335_
rlabel metal2 4200 17640 4200 17640 0 _0336_
rlabel metal2 46760 5600 46760 5600 0 _0337_
rlabel metal2 50456 4200 50456 4200 0 _0338_
rlabel metal2 57064 6160 57064 6160 0 _0339_
rlabel metal2 8568 22456 8568 22456 0 _0340_
rlabel metal2 8120 22736 8120 22736 0 _0341_
rlabel metal2 53704 8904 53704 8904 0 _0342_
rlabel metal2 19208 26152 19208 26152 0 _0343_
rlabel metal2 21952 12936 21952 12936 0 _0344_
rlabel metal2 52024 10920 52024 10920 0 _0345_
rlabel metal2 3528 21336 3528 21336 0 _0346_
rlabel metal2 50344 6160 50344 6160 0 _0347_
rlabel metal2 50792 6384 50792 6384 0 _0348_
rlabel metal2 51352 6328 51352 6328 0 _0349_
rlabel metal2 57176 7168 57176 7168 0 _0350_
rlabel metal3 57736 5096 57736 5096 0 _0351_
rlabel metal2 47096 5600 47096 5600 0 _0352_
rlabel metal2 47656 4760 47656 4760 0 _0353_
rlabel metal2 13384 24304 13384 24304 0 _0354_
rlabel metal3 48104 5880 48104 5880 0 _0355_
rlabel metal2 51128 6720 51128 6720 0 _0356_
rlabel metal2 53928 6104 53928 6104 0 _0357_
rlabel metal2 52248 5376 52248 5376 0 _0358_
rlabel metal2 52920 8624 52920 8624 0 _0359_
rlabel metal3 54880 10360 54880 10360 0 _0360_
rlabel metal3 21560 11368 21560 11368 0 _0361_
rlabel metal2 55272 5712 55272 5712 0 _0362_
rlabel metal2 57624 5824 57624 5824 0 _0363_
rlabel metal2 57848 3528 57848 3528 0 _0364_
rlabel metal2 18536 24080 18536 24080 0 _0365_
rlabel metal2 57960 3864 57960 3864 0 _0366_
rlabel metal2 55720 5936 55720 5936 0 _0367_
rlabel metal2 56168 6384 56168 6384 0 _0368_
rlabel metal2 54040 7112 54040 7112 0 _0369_
rlabel metal2 56504 8680 56504 8680 0 _0370_
rlabel metal2 48104 8120 48104 8120 0 _0371_
rlabel metal2 58184 7112 58184 7112 0 _0372_
rlabel metal2 56560 9800 56560 9800 0 _0373_
rlabel metal2 56392 10864 56392 10864 0 _0374_
rlabel metal3 56168 9688 56168 9688 0 _0375_
rlabel metal2 26264 23128 26264 23128 0 _0376_
rlabel metal2 48440 9688 48440 9688 0 _0377_
rlabel metal2 48552 8232 48552 8232 0 _0378_
rlabel metal2 48104 9968 48104 9968 0 _0379_
rlabel metal2 49560 9744 49560 9744 0 _0380_
rlabel metal2 21336 8624 21336 8624 0 _0381_
rlabel metal2 10696 8456 10696 8456 0 _0382_
rlabel metal2 9464 7952 9464 7952 0 _0383_
rlabel metal3 10136 8232 10136 8232 0 _0384_
rlabel metal2 10360 7896 10360 7896 0 _0385_
rlabel metal2 10472 5992 10472 5992 0 _0386_
rlabel metal2 2968 20496 2968 20496 0 _0387_
rlabel metal2 4088 7728 4088 7728 0 _0388_
rlabel metal2 3864 7840 3864 7840 0 _0389_
rlabel metal3 5320 7448 5320 7448 0 _0390_
rlabel metal2 6552 7504 6552 7504 0 _0391_
rlabel metal2 7784 7000 7784 7000 0 _0392_
rlabel metal2 10696 5824 10696 5824 0 _0393_
rlabel metal2 13160 3864 13160 3864 0 _0394_
rlabel metal3 13272 9912 13272 9912 0 _0395_
rlabel metal2 15960 6888 15960 6888 0 _0396_
rlabel metal2 12936 7560 12936 7560 0 _0397_
rlabel metal2 4760 20720 4760 20720 0 _0398_
rlabel metal2 12264 7392 12264 7392 0 _0399_
rlabel metal2 13608 5152 13608 5152 0 _0400_
rlabel metal3 9632 5096 9632 5096 0 _0401_
rlabel metal2 7616 6664 7616 6664 0 _0402_
rlabel metal2 6216 5824 6216 5824 0 _0403_
rlabel metal3 4200 5096 4200 5096 0 _0404_
rlabel metal2 5320 4816 5320 4816 0 _0405_
rlabel metal2 10248 5544 10248 5544 0 _0406_
rlabel metal3 5544 4312 5544 4312 0 _0407_
rlabel metal2 6664 4760 6664 4760 0 _0408_
rlabel metal2 2184 19376 2184 19376 0 _0409_
rlabel metal2 9016 5096 9016 5096 0 _0410_
rlabel metal3 11704 5376 11704 5376 0 _0411_
rlabel metal2 23688 8736 23688 8736 0 _0412_
rlabel metal2 4480 16296 4480 16296 0 _0413_
rlabel metal2 21112 15652 21112 15652 0 _0414_
rlabel metal2 4536 15484 4536 15484 0 _0415_
rlabel metal2 4312 14224 4312 14224 0 _0416_
rlabel metal2 4424 13720 4424 13720 0 _0417_
rlabel metal2 5096 13608 5096 13608 0 _0418_
rlabel metal2 18312 11480 18312 11480 0 _0419_
rlabel metal2 4648 20440 4648 20440 0 _0420_
rlabel metal3 21840 9128 21840 9128 0 _0421_
rlabel metal2 24472 9464 24472 9464 0 _0422_
rlabel metal2 8232 13608 8232 13608 0 _0423_
rlabel metal2 7000 15204 7000 15204 0 _0424_
rlabel metal2 8344 12880 8344 12880 0 _0425_
rlabel metal3 20832 10696 20832 10696 0 _0426_
rlabel metal2 9576 14168 9576 14168 0 _0427_
rlabel metal2 9128 13720 9128 13720 0 _0428_
rlabel metal2 21448 13216 21448 13216 0 _0429_
rlabel metal2 23016 11144 23016 11144 0 _0430_
rlabel metal2 8008 16744 8008 16744 0 _0431_
rlabel metal2 24136 8120 24136 8120 0 _0432_
rlabel metal2 23464 11256 23464 11256 0 _0433_
rlabel metal2 23352 11760 23352 11760 0 _0434_
rlabel metal2 24248 9408 24248 9408 0 _0435_
rlabel metal2 22008 9856 22008 9856 0 _0436_
rlabel metal2 25032 6720 25032 6720 0 _0437_
rlabel metal2 25928 8736 25928 8736 0 _0438_
rlabel metal2 26096 7448 26096 7448 0 _0439_
rlabel metal2 25816 7840 25816 7840 0 _0440_
rlabel metal3 26348 9128 26348 9128 0 _0441_
rlabel metal2 10360 20776 10360 20776 0 _0442_
rlabel metal3 26152 8904 26152 8904 0 _0443_
rlabel metal2 25144 5432 25144 5432 0 _0444_
rlabel metal2 23352 5768 23352 5768 0 _0445_
rlabel metal3 21504 5880 21504 5880 0 _0446_
rlabel metal2 25480 4760 25480 4760 0 _0447_
rlabel metal2 13944 10136 13944 10136 0 _0448_
rlabel metal2 15512 8344 15512 8344 0 _0449_
rlabel metal2 15288 7392 15288 7392 0 _0450_
rlabel metal3 16968 10360 16968 10360 0 _0451_
rlabel metal2 18088 10080 18088 10080 0 _0452_
rlabel metal2 17080 19600 17080 19600 0 _0453_
rlabel metal2 18144 7448 18144 7448 0 _0454_
rlabel metal2 15400 7728 15400 7728 0 _0455_
rlabel metal3 17864 6776 17864 6776 0 _0456_
rlabel metal2 16184 5656 16184 5656 0 _0457_
rlabel metal3 13160 4536 13160 4536 0 _0458_
rlabel metal2 13272 3976 13272 3976 0 _0459_
rlabel metal3 12936 4312 12936 4312 0 _0460_
rlabel metal2 10584 5488 10584 5488 0 _0461_
rlabel metal3 17304 4984 17304 4984 0 _0462_
rlabel metal2 6888 4032 6888 4032 0 _0463_
rlabel metal3 4872 18536 4872 18536 0 _0464_
rlabel metal2 8232 5544 8232 5544 0 _0465_
rlabel metal2 8008 5208 8008 5208 0 _0466_
rlabel metal3 15764 5096 15764 5096 0 _0467_
rlabel metal2 25256 4592 25256 4592 0 _0468_
rlabel metal2 24136 4200 24136 4200 0 _0469_
rlabel metal2 22120 5208 22120 5208 0 _0470_
rlabel metal2 18928 9016 18928 9016 0 _0471_
rlabel metal3 4704 9128 4704 9128 0 _0472_
rlabel metal2 4424 8904 4424 8904 0 _0473_
rlabel metal2 18312 8736 18312 8736 0 _0474_
rlabel metal2 1960 19040 1960 19040 0 _0475_
rlabel metal2 20552 5936 20552 5936 0 _0476_
rlabel metal2 21504 4424 21504 4424 0 _0477_
rlabel metal3 17248 4424 17248 4424 0 _0478_
rlabel metal3 20496 3752 20496 3752 0 _0479_
rlabel metal3 23128 4312 23128 4312 0 _0480_
rlabel metal2 18256 5992 18256 5992 0 _0481_
rlabel metal2 18816 5320 18816 5320 0 _0482_
rlabel metal2 17864 8176 17864 8176 0 _0483_
rlabel metal3 18704 5880 18704 5880 0 _0484_
rlabel metal2 19432 6104 19432 6104 0 _0485_
rlabel metal2 17920 18312 17920 18312 0 _0486_
rlabel metal2 19544 4816 19544 4816 0 _0487_
rlabel metal2 19992 4592 19992 4592 0 _0488_
rlabel metal2 20664 4984 20664 4984 0 _0489_
rlabel metal3 24752 4424 24752 4424 0 _0490_
rlabel metal3 22232 4088 22232 4088 0 _0491_
rlabel metal3 25144 4088 25144 4088 0 _0492_
rlabel metal2 26824 4256 26824 4256 0 _0493_
rlabel metal3 24808 3416 24808 3416 0 _0494_
rlabel metal2 25032 3528 25032 3528 0 _0495_
rlabel metal2 27384 3864 27384 3864 0 _0496_
rlabel metal2 16520 18816 16520 18816 0 _0497_
rlabel metal3 29456 7448 29456 7448 0 _0498_
rlabel metal2 25704 5040 25704 5040 0 _0499_
rlabel metal2 26040 5488 26040 5488 0 _0500_
rlabel metal2 28168 7112 28168 7112 0 _0501_
rlabel metal2 30632 5320 30632 5320 0 _0502_
rlabel metal3 32704 4312 32704 4312 0 _0503_
rlabel metal2 32984 3808 32984 3808 0 _0504_
rlabel metal2 33320 5712 33320 5712 0 _0505_
rlabel metal2 32480 5880 32480 5880 0 _0506_
rlabel metal3 34048 5656 34048 5656 0 _0507_
rlabel metal2 17584 23016 17584 23016 0 _0508_
rlabel metal2 27552 8120 27552 8120 0 _0509_
rlabel metal3 28448 8232 28448 8232 0 _0510_
rlabel metal2 28896 8120 28896 8120 0 _0511_
rlabel metal2 31976 6272 31976 6272 0 _0512_
rlabel metal2 31192 8176 31192 8176 0 _0513_
rlabel metal2 31080 8288 31080 8288 0 _0514_
rlabel metal2 31752 6328 31752 6328 0 _0515_
rlabel metal2 32816 5656 32816 5656 0 _0516_
rlabel metal2 33432 5432 33432 5432 0 _0517_
rlabel metal2 34944 5208 34944 5208 0 _0518_
rlabel metal3 7952 16856 7952 16856 0 _0519_
rlabel metal3 34944 7560 34944 7560 0 _0520_
rlabel metal2 34552 7728 34552 7728 0 _0521_
rlabel metal3 33488 7448 33488 7448 0 _0522_
rlabel metal2 33096 6944 33096 6944 0 _0523_
rlabel metal2 35224 7168 35224 7168 0 _0524_
rlabel metal2 49000 4704 49000 4704 0 _0525_
rlabel metal2 49336 10416 49336 10416 0 _0526_
rlabel metal2 50008 11424 50008 11424 0 _0527_
rlabel metal2 49336 9912 49336 9912 0 _0528_
rlabel metal2 53368 19264 53368 19264 0 _0529_
rlabel metal2 15288 22400 15288 22400 0 _0530_
rlabel metal2 55832 23576 55832 23576 0 _0531_
rlabel metal2 53704 25760 53704 25760 0 _0532_
rlabel metal2 54936 25256 54936 25256 0 _0533_
rlabel metal2 56784 23912 56784 23912 0 _0534_
rlabel metal2 56840 22176 56840 22176 0 _0535_
rlabel metal2 57176 23912 57176 23912 0 _0536_
rlabel metal2 53816 22288 53816 22288 0 _0537_
rlabel metal2 46536 22512 46536 22512 0 _0538_
rlabel metal2 48104 22680 48104 22680 0 _0539_
rlabel metal2 45080 19656 45080 19656 0 _0540_
rlabel metal2 17864 22456 17864 22456 0 _0541_
rlabel metal2 49056 20664 49056 20664 0 _0542_
rlabel metal2 47656 21616 47656 21616 0 _0543_
rlabel metal2 51632 20776 51632 20776 0 _0544_
rlabel metal2 52808 17696 52808 17696 0 _0545_
rlabel metal2 44744 18088 44744 18088 0 _0546_
rlabel metal2 47320 22680 47320 22680 0 _0547_
rlabel metal2 47096 23464 47096 23464 0 _0548_
rlabel metal2 49224 18368 49224 18368 0 _0549_
rlabel metal2 45640 18088 45640 18088 0 _0550_
rlabel metal2 46984 22792 46984 22792 0 _0551_
rlabel metal2 22680 20216 22680 20216 0 _0552_
rlabel metal2 45528 18928 45528 18928 0 _0553_
rlabel via2 42840 18536 42840 18536 0 _0554_
rlabel metal3 44856 18424 44856 18424 0 _0555_
rlabel metal2 45192 17416 45192 17416 0 _0556_
rlabel metal2 43512 16968 43512 16968 0 _0557_
rlabel metal2 42504 16912 42504 16912 0 _0558_
rlabel metal2 42616 17472 42616 17472 0 _0559_
rlabel metal2 43960 16408 43960 16408 0 _0560_
rlabel metal2 49336 16016 49336 16016 0 _0561_
rlabel metal2 49448 18032 49448 18032 0 _0562_
rlabel metal2 29736 22624 29736 22624 0 _0563_
rlabel metal2 47208 18424 47208 18424 0 _0564_
rlabel metal2 47824 16744 47824 16744 0 _0565_
rlabel metal3 48832 20104 48832 20104 0 _0566_
rlabel metal2 48104 17360 48104 17360 0 _0567_
rlabel metal2 47880 15736 47880 15736 0 _0568_
rlabel metal2 47768 21056 47768 21056 0 _0569_
rlabel metal2 48104 19096 48104 19096 0 _0570_
rlabel metal2 50568 18704 50568 18704 0 _0571_
rlabel metal2 49000 15680 49000 15680 0 _0572_
rlabel metal2 53368 18200 53368 18200 0 _0573_
rlabel metal2 3192 9688 3192 9688 0 _0574_
rlabel metal2 53928 19320 53928 19320 0 _0575_
rlabel metal2 54040 20440 54040 20440 0 _0576_
rlabel metal2 54152 25368 54152 25368 0 _0577_
rlabel metal2 55440 22232 55440 22232 0 _0578_
rlabel metal2 56504 21504 56504 21504 0 _0579_
rlabel metal2 55720 20720 55720 20720 0 _0580_
rlabel metal2 57064 17136 57064 17136 0 _0581_
rlabel metal2 57960 21168 57960 21168 0 _0582_
rlabel metal2 57288 22232 57288 22232 0 _0583_
rlabel metal2 58128 19208 58128 19208 0 _0584_
rlabel metal2 3304 7168 3304 7168 0 _0585_
rlabel metal2 57568 19096 57568 19096 0 _0586_
rlabel metal2 55832 17192 55832 17192 0 _0587_
rlabel metal2 54376 21336 54376 21336 0 _0588_
rlabel metal2 54040 22008 54040 22008 0 _0589_
rlabel metal2 53760 15288 53760 15288 0 _0590_
rlabel metal2 55496 21616 55496 21616 0 _0591_
rlabel metal3 56280 16744 56280 16744 0 _0592_
rlabel metal2 53480 15736 53480 15736 0 _0593_
rlabel metal2 54600 17752 54600 17752 0 _0594_
rlabel metal2 53144 18536 53144 18536 0 _0595_
rlabel metal2 2520 7896 2520 7896 0 _0596_
rlabel metal2 53480 20104 53480 20104 0 _0597_
rlabel metal2 54936 16856 54936 16856 0 _0598_
rlabel metal2 54712 15792 54712 15792 0 _0599_
rlabel metal2 55384 16352 55384 16352 0 _0600_
rlabel metal2 49896 13888 49896 13888 0 _0601_
rlabel metal2 55048 14616 55048 14616 0 _0602_
rlabel metal2 55048 13216 55048 13216 0 _0603_
rlabel metal3 56896 14504 56896 14504 0 _0604_
rlabel metal2 55328 15848 55328 15848 0 _0605_
rlabel metal2 48776 13944 48776 13944 0 _0606_
rlabel metal3 18648 9912 18648 9912 0 _0607_
rlabel metal2 49224 15232 49224 15232 0 _0608_
rlabel metal2 48776 15148 48776 15148 0 _0609_
rlabel metal2 48888 12432 48888 12432 0 _0610_
rlabel metal2 49168 9800 49168 9800 0 _0611_
rlabel metal2 55048 16912 55048 16912 0 _0612_
rlabel metal3 45416 8176 45416 8176 0 _0613_
rlabel metal2 55832 13440 55832 13440 0 _0614_
rlabel metal3 56728 12264 56728 12264 0 _0615_
rlabel metal3 56392 12152 56392 12152 0 _0616_
rlabel metal3 15400 13552 15400 13552 0 _0617_
rlabel metal2 35672 6384 35672 6384 0 _0618_
rlabel metal2 45528 10416 45528 10416 0 _0619_
rlabel metal2 58184 12096 58184 12096 0 _0620_
rlabel metal3 56448 11144 56448 11144 0 _0621_
rlabel metal2 57736 16044 57736 16044 0 _0622_
rlabel metal3 57232 16856 57232 16856 0 _0623_
rlabel metal2 33600 8344 33600 8344 0 _0624_
rlabel metal3 55888 17080 55888 17080 0 _0625_
rlabel metal3 16968 23016 16968 23016 0 _0626_
rlabel metal2 56056 11760 56056 11760 0 _0627_
rlabel metal2 55832 11284 55832 11284 0 _0628_
rlabel metal2 35896 9688 35896 9688 0 _0629_
rlabel metal2 55608 11424 55608 11424 0 _0630_
rlabel metal2 57288 11928 57288 11928 0 _0631_
rlabel metal2 52864 13048 52864 13048 0 _0632_
rlabel metal2 35784 5600 35784 5600 0 _0633_
rlabel metal2 45416 6272 45416 6272 0 _0634_
rlabel metal3 55608 12824 55608 12824 0 _0635_
rlabel metal2 10248 18592 10248 18592 0 _0636_
rlabel metal2 29736 5992 29736 5992 0 _0637_
rlabel metal2 29064 4480 29064 4480 0 _0638_
rlabel metal2 49896 4704 49896 4704 0 _0639_
rlabel metal2 45304 7840 45304 7840 0 _0640_
rlabel metal2 42560 9800 42560 9800 0 _0641_
rlabel metal3 44184 7560 44184 7560 0 _0642_
rlabel metal2 45416 7672 45416 7672 0 _0643_
rlabel metal2 46424 7952 46424 7952 0 _0644_
rlabel metal2 45976 8568 45976 8568 0 _0645_
rlabel metal2 18928 11480 18928 11480 0 _0646_
rlabel metal2 49000 9072 49000 9072 0 _0647_
rlabel metal2 41440 17640 41440 17640 0 _0648_
rlabel metal2 43736 16408 43736 16408 0 _0649_
rlabel metal2 45752 15624 45752 15624 0 _0650_
rlabel metal2 45864 14728 45864 14728 0 _0651_
rlabel metal2 48776 9576 48776 9576 0 _0652_
rlabel metal2 49392 5208 49392 5208 0 _0653_
rlabel metal2 27832 4984 27832 4984 0 _0654_
rlabel metal2 48888 5600 48888 5600 0 _0655_
rlabel metal2 16408 15568 16408 15568 0 _0656_
rlabel metal2 44296 7168 44296 7168 0 _0657_
rlabel metal2 46760 7448 46760 7448 0 _0658_
rlabel metal2 47208 7952 47208 7952 0 _0659_
rlabel metal3 48608 8232 48608 8232 0 _0660_
rlabel metal2 48272 15960 48272 15960 0 _0661_
rlabel metal2 49112 8456 49112 8456 0 _0662_
rlabel metal2 49224 6384 49224 6384 0 _0663_
rlabel metal3 15904 15400 15904 15400 0 _0664_
rlabel metal2 15960 21112 15960 21112 0 _0665_
rlabel metal2 15008 22120 15008 22120 0 _0666_
rlabel metal2 18424 24136 18424 24136 0 _0667_
rlabel metal2 17528 25480 17528 25480 0 _0668_
rlabel metal2 15736 24192 15736 24192 0 _0669_
rlabel metal2 22456 23744 22456 23744 0 _0670_
rlabel metal2 3080 16352 3080 16352 0 _0671_
rlabel metal2 2352 8120 2352 8120 0 _0672_
rlabel metal3 19208 12096 19208 12096 0 _0673_
rlabel metal2 19880 8456 19880 8456 0 _0674_
rlabel metal2 20216 17808 20216 17808 0 _0675_
rlabel metal2 19768 24248 19768 24248 0 _0676_
rlabel metal2 17752 22568 17752 22568 0 _0677_
rlabel metal2 19096 25368 19096 25368 0 _0678_
rlabel metal3 23520 23800 23520 23800 0 _0679_
rlabel metal2 12376 24248 12376 24248 0 _0680_
rlabel metal2 10696 20328 10696 20328 0 _0681_
rlabel metal2 10136 20888 10136 20888 0 _0682_
rlabel metal2 11928 22848 11928 22848 0 _0683_
rlabel metal2 20664 18928 20664 18928 0 _0684_
rlabel metal3 9352 26264 9352 26264 0 _0685_
rlabel metal2 11816 21504 11816 21504 0 _0686_
rlabel metal2 11032 18032 11032 18032 0 _0687_
rlabel metal2 7112 17976 7112 17976 0 _0688_
rlabel metal2 8232 17752 8232 17752 0 _0689_
rlabel metal3 10080 17640 10080 17640 0 _0690_
rlabel metal2 11480 22512 11480 22512 0 _0691_
rlabel metal3 1246 1400 1246 1400 0 a[0]
rlabel metal3 1302 3192 1302 3192 0 a[1]
rlabel metal2 1848 4816 1848 4816 0 a[2]
rlabel metal3 1736 6720 1736 6720 0 a[3]
rlabel metal2 2744 8792 2744 8792 0 a[4]
rlabel metal2 1960 9744 1960 9744 0 a[5]
rlabel metal2 1960 12880 1960 12880 0 a[6]
rlabel metal2 1736 10864 1736 10864 0 a[7]
rlabel metal2 1680 15848 1680 15848 0 b[0]
rlabel metal2 1848 16240 1848 16240 0 b[1]
rlabel metal2 1736 19264 1736 19264 0 b[2]
rlabel metal3 1302 21112 1302 21112 0 b[3]
rlabel metal2 2576 24696 2576 24696 0 b[4]
rlabel metal2 1736 25088 1736 25088 0 b[5]
rlabel metal2 2184 24864 2184 24864 0 b[6]
rlabel metal3 3150 28280 3150 28280 0 b[7]
rlabel metal2 3080 9184 3080 9184 0 net1
rlabel metal2 3192 17080 3192 17080 0 net10
rlabel metal2 2240 17864 2240 17864 0 net11
rlabel metal2 2296 16520 2296 16520 0 net12
rlabel metal2 1736 23856 1736 23856 0 net13
rlabel metal2 2744 16576 2744 16576 0 net14
rlabel metal2 2520 16464 2520 16464 0 net15
rlabel metal2 1288 19600 1288 19600 0 net16
rlabel metal2 47656 25928 47656 25928 0 net17
rlabel metal3 43568 26152 43568 26152 0 net18
rlabel metal2 50680 25536 50680 25536 0 net19
rlabel metal2 2072 5264 2072 5264 0 net2
rlabel metal2 55664 3528 55664 3528 0 net20
rlabel metal3 52976 5880 52976 5880 0 net21
rlabel metal2 49672 10304 49672 10304 0 net22
rlabel metal2 57624 13048 57624 13048 0 net23
rlabel metal2 57176 15960 57176 15960 0 net24
rlabel metal2 56672 19992 56672 19992 0 net25
rlabel metal2 54483 16520 54483 16520 0 net26
rlabel metal2 46480 18200 46480 18200 0 net27
rlabel metal2 17192 16296 17192 16296 0 net28
rlabel metal2 30576 25480 30576 25480 0 net29
rlabel metal2 15288 12096 15288 12096 0 net3
rlabel metal2 13272 25928 13272 25928 0 net30
rlabel metal3 7616 23128 7616 23128 0 net31
rlabel metal3 15148 24696 15148 24696 0 net32
rlabel metal2 49448 19544 49448 19544 0 net33
rlabel metal2 43624 21952 43624 21952 0 net34
rlabel metal2 15848 17864 15848 17864 0 net35
rlabel metal2 18312 23072 18312 23072 0 net36
rlabel metal2 20888 21840 20888 21840 0 net37
rlabel metal2 21560 16016 21560 16016 0 net38
rlabel metal3 21504 15960 21504 15960 0 net39
rlabel metal2 2296 23408 2296 23408 0 net4
rlabel metal3 16968 13944 16968 13944 0 net40
rlabel metal2 16128 14504 16128 14504 0 net41
rlabel metal2 23912 24640 23912 24640 0 net42
rlabel metal3 41160 19992 41160 19992 0 net43
rlabel metal2 48664 23856 48664 23856 0 net44
rlabel metal2 21112 24584 21112 24584 0 net45
rlabel metal2 38920 25816 38920 25816 0 net46
rlabel metal3 23184 21448 23184 21448 0 net47
rlabel metal2 27272 25144 27272 25144 0 net48
rlabel metal2 12936 25088 12936 25088 0 net49
rlabel metal2 1848 19432 1848 19432 0 net5
rlabel metal2 10808 23184 10808 23184 0 net50
rlabel metal2 2520 9184 2520 9184 0 net6
rlabel metal2 2744 13496 2744 13496 0 net7
rlabel metal2 2296 14224 2296 14224 0 net8
rlabel metal3 2464 15400 2464 15400 0 net9
rlabel metal2 1512 19712 1512 19712 0 op[0]
rlabel metal2 29848 28070 29848 28070 0 op[1]
rlabel metal2 50064 27272 50064 27272 0 op[2]
rlabel metal3 59234 2296 59234 2296 0 out[0]
rlabel metal3 58674 5880 58674 5880 0 out[1]
rlabel metal2 57960 10248 57960 10248 0 out[2]
rlabel metal2 57288 13384 57288 13384 0 out[3]
rlabel metal2 58072 16016 58072 16016 0 out[4]
rlabel metal3 57736 20160 57736 20160 0 out[5]
rlabel metal3 58450 23800 58450 23800 0 out[6]
rlabel metal3 58506 27384 58506 27384 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 60000 30000
<< end >>
