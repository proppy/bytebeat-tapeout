VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpu8_wrap
  CLASS BLOCK ;
  FOREIGN fpu8_wrap ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 150.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 4.000 7.280 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 4.000 16.240 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 4.000 25.200 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.440 4.000 70.000 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 4.000 96.880 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END b[7]
  PIN op[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 146.000 49.840 150.000 ;
    END
  END op[0]
  PIN op[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 146.000 149.520 150.000 ;
    END
  END op[1]
  PIN op[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 146.000 249.200 150.000 ;
    END
  END op[2]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 11.200 300.000 11.760 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 29.120 300.000 29.680 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 47.040 300.000 47.600 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 64.960 300.000 65.520 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 82.880 300.000 83.440 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 100.800 300.000 101.360 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 118.720 300.000 119.280 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 136.640 300.000 137.200 ;
    END
  END out[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 41.685 15.380 43.285 133.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 113.220 15.380 114.820 133.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.755 15.380 186.355 133.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 256.290 15.380 257.890 133.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 77.450 15.380 79.050 133.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 148.985 15.380 150.585 133.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 220.520 15.380 222.120 133.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 292.055 15.380 293.655 133.580 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 293.655 134.250 ;
      LAYER Metal2 ;
        RECT 6.300 145.700 48.980 146.000 ;
        RECT 50.140 145.700 148.660 146.000 ;
        RECT 149.820 145.700 248.340 146.000 ;
        RECT 249.500 145.700 293.515 146.000 ;
        RECT 6.300 6.810 293.515 145.700 ;
      LAYER Metal3 ;
        RECT 4.300 140.820 296.660 141.540 ;
        RECT 4.000 137.500 296.660 140.820 ;
        RECT 4.000 136.340 295.700 137.500 ;
        RECT 4.000 133.020 296.660 136.340 ;
        RECT 4.300 131.860 296.660 133.020 ;
        RECT 4.000 124.060 296.660 131.860 ;
        RECT 4.300 122.900 296.660 124.060 ;
        RECT 4.000 119.580 296.660 122.900 ;
        RECT 4.000 118.420 295.700 119.580 ;
        RECT 4.000 115.100 296.660 118.420 ;
        RECT 4.300 113.940 296.660 115.100 ;
        RECT 4.000 106.140 296.660 113.940 ;
        RECT 4.300 104.980 296.660 106.140 ;
        RECT 4.000 101.660 296.660 104.980 ;
        RECT 4.000 100.500 295.700 101.660 ;
        RECT 4.000 97.180 296.660 100.500 ;
        RECT 4.300 96.020 296.660 97.180 ;
        RECT 4.000 88.220 296.660 96.020 ;
        RECT 4.300 87.060 296.660 88.220 ;
        RECT 4.000 83.740 296.660 87.060 ;
        RECT 4.000 82.580 295.700 83.740 ;
        RECT 4.000 79.260 296.660 82.580 ;
        RECT 4.300 78.100 296.660 79.260 ;
        RECT 4.000 70.300 296.660 78.100 ;
        RECT 4.300 69.140 296.660 70.300 ;
        RECT 4.000 65.820 296.660 69.140 ;
        RECT 4.000 64.660 295.700 65.820 ;
        RECT 4.000 61.340 296.660 64.660 ;
        RECT 4.300 60.180 296.660 61.340 ;
        RECT 4.000 52.380 296.660 60.180 ;
        RECT 4.300 51.220 296.660 52.380 ;
        RECT 4.000 47.900 296.660 51.220 ;
        RECT 4.000 46.740 295.700 47.900 ;
        RECT 4.000 43.420 296.660 46.740 ;
        RECT 4.300 42.260 296.660 43.420 ;
        RECT 4.000 34.460 296.660 42.260 ;
        RECT 4.300 33.300 296.660 34.460 ;
        RECT 4.000 29.980 296.660 33.300 ;
        RECT 4.000 28.820 295.700 29.980 ;
        RECT 4.000 25.500 296.660 28.820 ;
        RECT 4.300 24.340 296.660 25.500 ;
        RECT 4.000 16.540 296.660 24.340 ;
        RECT 4.300 15.380 296.660 16.540 ;
        RECT 4.000 12.060 296.660 15.380 ;
        RECT 4.000 10.900 295.700 12.060 ;
        RECT 4.000 7.580 296.660 10.900 ;
        RECT 4.300 6.860 296.660 7.580 ;
      LAYER Metal4 ;
        RECT 9.100 26.970 41.385 131.510 ;
        RECT 43.585 26.970 77.150 131.510 ;
        RECT 79.350 26.970 112.920 131.510 ;
        RECT 115.120 26.970 148.685 131.510 ;
        RECT 150.885 26.970 184.455 131.510 ;
        RECT 186.655 26.970 220.220 131.510 ;
        RECT 222.420 26.970 255.990 131.510 ;
        RECT 258.190 26.970 279.860 131.510 ;
  END
END fpu8_wrap
END LIBRARY

